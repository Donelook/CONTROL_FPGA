-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 5 2025 21:16:21

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T45 : out std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    T01 : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__45224\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44951\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44939\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44855\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44380\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44290\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44110\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44107\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43535\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43307\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43214\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43049\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42668\ : std_logic;
signal \N__42665\ : std_logic;
signal \N__42662\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42457\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41906\ : std_logic;
signal \N__41903\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41681\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38746\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \N_38_i_i\ : std_logic;
signal \rgb_drv_RNOZ0\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_3_10_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_3_11_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_154\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_149\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_153\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_53\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_155\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI3VBED1_0_16_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIP1MD11_0_12_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIP1MD11_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNINVLD11_0_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIQ2MD11_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNI51CED1_0_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_\ : std_logic;
signal \bfn_7_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_f0_i_1Z0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNINVLD11_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_315\ : std_logic;
signal \elapsed_time_ns_1_RNIO0MD11_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIR4ND11_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNIS5ND11_0_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14\ : std_logic;
signal \elapsed_time_ns_1_RNI1TBED1_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI1TBED1_0_14_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIL13KD1_0_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal s4_phy_c : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \elapsed_time_ns_1_RNI40CED1_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI51CED1_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI3VBED1_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3Z0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_328\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \elapsed_time_ns_1_RNI1BND11_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNIP2ND11_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNI1BND11_0_29_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_o5_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_o5_7Z0Z_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \elapsed_time_ns_1_RNIO1ND11_0_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \elapsed_time_ns_1_RNIQ3ND11_0_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \elapsed_time_ns_1_RNIT6ND11_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNIT6ND11_0_25_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_o5_6Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \elapsed_time_ns_1_RNIV8ND11_0_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \elapsed_time_ns_1_RNIU7ND11_0_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \elapsed_time_ns_1_RNI0AND11_0_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \elapsed_time_ns_1_RNIP3OD11_0_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_432_i_g\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_432_i\ : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal s3_phy_c : std_logic;
signal il_min_comp1_c : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \elapsed_time_ns_1_RNI62CED1_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a5_1_1_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_325_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNIS4MD11_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_307_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_45_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \T12_c\ : std_logic;
signal state_ns_i_a3_1 : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_stoper_state12_1_0_i\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \elapsed_time_ns_1_RNID6DJ11_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNID6DJ11_0_7_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\ : std_logic;
signal \elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_i_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNIA3DJ11_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \elapsed_time_ns_1_RNIB4DJ11_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \elapsed_time_ns_1_RNIE7DJ11_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \elapsed_time_ns_1_RNIQ4OD11_0_31\ : std_logic;
signal \elapsed_time_ns_1_RNIDP2KD1_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_f0_0_1Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_325\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_327\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_7_f0_0_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_433_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \elapsed_time_ns_1_RNI81DJ11_0_2\ : std_logic;
signal \elapsed_time_ns_1_RNI81DJ11_0_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIQURR91_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_283\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst1.N_56\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_RNOZ0Z_0_cascade_\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_0_sqmuxa_cascade_\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_7\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_9\ : std_logic;
signal start_stop_c : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal \T23_c\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74_16_cascade_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHEZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18\ : std_logic;
signal \current_shift_inst.control_input_1_axb_0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19\ : std_logic;
signal \current_shift_inst.control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20\ : std_logic;
signal \current_shift_inst.control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22\ : std_logic;
signal \current_shift_inst.control_input_1_axb_3\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23\ : std_logic;
signal \current_shift_inst.control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24\ : std_logic;
signal \current_shift_inst.control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26\ : std_logic;
signal \current_shift_inst.control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27\ : std_logic;
signal \current_shift_inst.control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_30\ : std_logic;
signal \phase_controller_inst2.time_passed_RNI9M3O\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \T01_c\ : std_logic;
signal s1_phy_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \T45_c\ : std_logic;
signal \current_shift_inst.timer_s1.N_166_i\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_62\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_72\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_31\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_45\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal state_3 : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_13_27_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_167_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_358_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\ : std_logic;
signal \elapsed_time_ns_1_RNIFJ2591_0_7_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_382_i\ : std_logic;
signal \elapsed_time_ns_1_RNIIU2KD1_0_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_235_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_stoper_state12_1_0_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.N_45\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_219\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_12\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_23\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_0_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_30\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_363_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI3JIF91_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNIRBJF91_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNIRAIF91_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNI3JIF91_0_29_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIQ9IF91_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNISBIF91_0_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_o5_7Z0Z_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_381\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_359_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_381_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_251_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIDH2591_0_5_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_241_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIPFL2M1_0_1\ : std_logic;
signal \elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_f0_0_1Z0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_103\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_380\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_341\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_367\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_367_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_378\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_349\ : std_logic;
signal \elapsed_time_ns_1_RNIVEIF91_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_o5_6Z0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNI2IIF91_0_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_345\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_348\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_347\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_347_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_365\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNI0GIF91_0_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNITCIF91_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNI1HIF91_0_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNIUDIF91_0_24\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_434_i\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.N_55\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\ : std_logic;
signal \elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI1OL2M1_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_244\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_249_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIFJ2591_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNIGK2591_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIUKL2M1_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_250\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_f0_i_1Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9\ : std_logic;
signal \elapsed_time_ns_1_RNIAE2591_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2\ : std_logic;
signal \elapsed_time_ns_1_RNIRHL2M1_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIUCHF91_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNIDH2591_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_249\ : std_logic;
signal \elapsed_time_ns_1_RNICG2591_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.N_166_i_g\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_434_i_g\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_stoper_state12_1_0_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.N_1310_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.N_45_cascade_\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_18_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_18_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_18_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_435_i\ : std_logic;
signal \elapsed_time_ns_1_RNIR9HF91_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNIDE4DM1_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNIP7HF91_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIQ8HF91_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIFG4DM1_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_241\ : std_logic;
signal \elapsed_time_ns_1_RNISAHF91_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNIIJ4DM1_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNIHI4DM1_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNIGH4DM1_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNISCJF91_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal red_c_g : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84ADZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_18_21_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_stoper_state12_1_0_i\ : std_logic;

signal reset_wire : std_logic;
signal \T01_wire\ : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal \T12_wire\ : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal \T45_wire\ : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal rgb_b_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    T01 <= \T01_wire\;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    T12 <= \T12_wire\;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    T45 <= \T45_wire\;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    rgb_b <= rgb_b_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__19364\&\N__19357\&\N__19362\&\N__19356\&\N__19363\&\N__19355\&\N__19365\&\N__19352\&\N__19358\&\N__19351\&\N__19359\&\N__19353\&\N__19360\&\N__19354\&\N__19361\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__40615\&\N__40611\&'0'&'0'&'0'&\N__40609\&\N__40614\&\N__40610\&\N__40613\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__19411\&\N__19416\&\N__19412\&\N__19417\&\N__19413\&\N__19782\&\N__19692\&\N__19737\&\N__19767\&\N__18231\&\N__19540\&\N__18813\&\N__19102\&\N__19117\&\N__19132\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__40468\&\N__40465\&'0'&'0'&'0'&\N__40463\&\N__40467\&\N__40464\&\N__40466\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__20453\,
            RESETB => \N__28073\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__40612\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__40608\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__40469\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__40462\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__45222\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45224\,
            DIN => \N__45223\,
            DOUT => \N__45222\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__45224\,
            PADOUT => \N__45223\,
            PADIN => \N__45222\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T01_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45213\,
            DIN => \N__45212\,
            DOUT => \N__45211\,
            PACKAGEPIN => \T01_wire\
        );

    \T01_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__45213\,
            PADOUT => \N__45212\,
            PADIN => \N__45211\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27986\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45204\,
            DIN => \N__45203\,
            DOUT => \N__45202\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__45204\,
            PADOUT => \N__45203\,
            PADIN => \N__45202\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45195\,
            DIN => \N__45194\,
            DOUT => \N__45193\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__45195\,
            PADOUT => \N__45194\,
            PADIN => \N__45193\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45186\,
            DIN => \N__45185\,
            DOUT => \N__45184\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__45186\,
            PADOUT => \N__45185\,
            PADIN => \N__45184\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26549\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45177\,
            DIN => \N__45176\,
            DOUT => \N__45175\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__45177\,
            PADOUT => \N__45176\,
            PADIN => \N__45175\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20345\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45168\,
            DIN => \N__45167\,
            DOUT => \N__45166\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__45168\,
            PADOUT => \N__45167\,
            PADIN => \N__45166\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45159\,
            DIN => \N__45158\,
            DOUT => \N__45157\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__45159\,
            PADOUT => \N__45158\,
            PADIN => \N__45157\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29384\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45150\,
            DIN => \N__45149\,
            DOUT => \N__45148\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__45150\,
            PADOUT => \N__45149\,
            PADIN => \N__45148\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25076\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45141\,
            DIN => \N__45140\,
            DOUT => \N__45139\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__45141\,
            PADOUT => \N__45140\,
            PADIN => \N__45139\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45132\,
            DIN => \N__45131\,
            DOUT => \N__45130\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__45132\,
            PADOUT => \N__45131\,
            PADIN => \N__45130\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27962\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45123\,
            DIN => \N__45122\,
            DOUT => \N__45121\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__45123\,
            PADOUT => \N__45122\,
            PADIN => \N__45121\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23114\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45114\,
            DIN => \N__45113\,
            DOUT => \N__45112\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__45114\,
            PADOUT => \N__45113\,
            PADIN => \N__45112\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45105\,
            DIN => \N__45104\,
            DOUT => \N__45103\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__45105\,
            PADOUT => \N__45104\,
            PADIN => \N__45103\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23906\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T45_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45096\,
            DIN => \N__45095\,
            DOUT => \N__45094\,
            PACKAGEPIN => \T45_wire\
        );

    \T45_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__45096\,
            PADOUT => \N__45095\,
            PADIN => \N__45094\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27854\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45087\,
            DIN => \N__45086\,
            DOUT => \N__45085\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__45087\,
            PADOUT => \N__45086\,
            PADIN => \N__45085\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__45078\,
            DIN => \N__45077\,
            DOUT => \N__45076\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__45078\,
            PADOUT => \N__45077\,
            PADIN => \N__45076\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__10663\ : InMux
    port map (
            O => \N__45059\,
            I => \N__45055\
        );

    \I__10662\ : InMux
    port map (
            O => \N__45058\,
            I => \N__45052\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__45055\,
            I => \N__45049\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__45052\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__10659\ : Odrv4
    port map (
            O => \N__45049\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__10658\ : InMux
    port map (
            O => \N__45044\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__10657\ : InMux
    port map (
            O => \N__45041\,
            I => \N__45037\
        );

    \I__10656\ : InMux
    port map (
            O => \N__45040\,
            I => \N__45034\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__45037\,
            I => \N__45031\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__45034\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__10653\ : Odrv12
    port map (
            O => \N__45031\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__10652\ : InMux
    port map (
            O => \N__45026\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__10651\ : InMux
    port map (
            O => \N__45023\,
            I => \N__45019\
        );

    \I__10650\ : InMux
    port map (
            O => \N__45022\,
            I => \N__45016\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__45019\,
            I => \N__45013\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__45016\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__10647\ : Odrv12
    port map (
            O => \N__45013\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__10646\ : InMux
    port map (
            O => \N__45008\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__10645\ : InMux
    port map (
            O => \N__45005\,
            I => \N__45001\
        );

    \I__10644\ : InMux
    port map (
            O => \N__45004\,
            I => \N__44998\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__45001\,
            I => \N__44995\
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__44998\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__10641\ : Odrv4
    port map (
            O => \N__44995\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__10640\ : InMux
    port map (
            O => \N__44990\,
            I => \bfn_18_21_0_\
        );

    \I__10639\ : InMux
    port map (
            O => \N__44987\,
            I => \N__44983\
        );

    \I__10638\ : InMux
    port map (
            O => \N__44986\,
            I => \N__44980\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__44983\,
            I => \N__44977\
        );

    \I__10636\ : LocalMux
    port map (
            O => \N__44980\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__44977\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10634\ : InMux
    port map (
            O => \N__44972\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__10633\ : InMux
    port map (
            O => \N__44969\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__10632\ : InMux
    port map (
            O => \N__44966\,
            I => \N__44962\
        );

    \I__10631\ : InMux
    port map (
            O => \N__44965\,
            I => \N__44959\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__44962\,
            I => \N__44956\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__44959\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10628\ : Odrv4
    port map (
            O => \N__44956\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10627\ : ClkMux
    port map (
            O => \N__44951\,
            I => \N__44591\
        );

    \I__10626\ : ClkMux
    port map (
            O => \N__44950\,
            I => \N__44591\
        );

    \I__10625\ : ClkMux
    port map (
            O => \N__44949\,
            I => \N__44591\
        );

    \I__10624\ : ClkMux
    port map (
            O => \N__44948\,
            I => \N__44591\
        );

    \I__10623\ : ClkMux
    port map (
            O => \N__44947\,
            I => \N__44591\
        );

    \I__10622\ : ClkMux
    port map (
            O => \N__44946\,
            I => \N__44591\
        );

    \I__10621\ : ClkMux
    port map (
            O => \N__44945\,
            I => \N__44591\
        );

    \I__10620\ : ClkMux
    port map (
            O => \N__44944\,
            I => \N__44591\
        );

    \I__10619\ : ClkMux
    port map (
            O => \N__44943\,
            I => \N__44591\
        );

    \I__10618\ : ClkMux
    port map (
            O => \N__44942\,
            I => \N__44591\
        );

    \I__10617\ : ClkMux
    port map (
            O => \N__44941\,
            I => \N__44591\
        );

    \I__10616\ : ClkMux
    port map (
            O => \N__44940\,
            I => \N__44591\
        );

    \I__10615\ : ClkMux
    port map (
            O => \N__44939\,
            I => \N__44591\
        );

    \I__10614\ : ClkMux
    port map (
            O => \N__44938\,
            I => \N__44591\
        );

    \I__10613\ : ClkMux
    port map (
            O => \N__44937\,
            I => \N__44591\
        );

    \I__10612\ : ClkMux
    port map (
            O => \N__44936\,
            I => \N__44591\
        );

    \I__10611\ : ClkMux
    port map (
            O => \N__44935\,
            I => \N__44591\
        );

    \I__10610\ : ClkMux
    port map (
            O => \N__44934\,
            I => \N__44591\
        );

    \I__10609\ : ClkMux
    port map (
            O => \N__44933\,
            I => \N__44591\
        );

    \I__10608\ : ClkMux
    port map (
            O => \N__44932\,
            I => \N__44591\
        );

    \I__10607\ : ClkMux
    port map (
            O => \N__44931\,
            I => \N__44591\
        );

    \I__10606\ : ClkMux
    port map (
            O => \N__44930\,
            I => \N__44591\
        );

    \I__10605\ : ClkMux
    port map (
            O => \N__44929\,
            I => \N__44591\
        );

    \I__10604\ : ClkMux
    port map (
            O => \N__44928\,
            I => \N__44591\
        );

    \I__10603\ : ClkMux
    port map (
            O => \N__44927\,
            I => \N__44591\
        );

    \I__10602\ : ClkMux
    port map (
            O => \N__44926\,
            I => \N__44591\
        );

    \I__10601\ : ClkMux
    port map (
            O => \N__44925\,
            I => \N__44591\
        );

    \I__10600\ : ClkMux
    port map (
            O => \N__44924\,
            I => \N__44591\
        );

    \I__10599\ : ClkMux
    port map (
            O => \N__44923\,
            I => \N__44591\
        );

    \I__10598\ : ClkMux
    port map (
            O => \N__44922\,
            I => \N__44591\
        );

    \I__10597\ : ClkMux
    port map (
            O => \N__44921\,
            I => \N__44591\
        );

    \I__10596\ : ClkMux
    port map (
            O => \N__44920\,
            I => \N__44591\
        );

    \I__10595\ : ClkMux
    port map (
            O => \N__44919\,
            I => \N__44591\
        );

    \I__10594\ : ClkMux
    port map (
            O => \N__44918\,
            I => \N__44591\
        );

    \I__10593\ : ClkMux
    port map (
            O => \N__44917\,
            I => \N__44591\
        );

    \I__10592\ : ClkMux
    port map (
            O => \N__44916\,
            I => \N__44591\
        );

    \I__10591\ : ClkMux
    port map (
            O => \N__44915\,
            I => \N__44591\
        );

    \I__10590\ : ClkMux
    port map (
            O => \N__44914\,
            I => \N__44591\
        );

    \I__10589\ : ClkMux
    port map (
            O => \N__44913\,
            I => \N__44591\
        );

    \I__10588\ : ClkMux
    port map (
            O => \N__44912\,
            I => \N__44591\
        );

    \I__10587\ : ClkMux
    port map (
            O => \N__44911\,
            I => \N__44591\
        );

    \I__10586\ : ClkMux
    port map (
            O => \N__44910\,
            I => \N__44591\
        );

    \I__10585\ : ClkMux
    port map (
            O => \N__44909\,
            I => \N__44591\
        );

    \I__10584\ : ClkMux
    port map (
            O => \N__44908\,
            I => \N__44591\
        );

    \I__10583\ : ClkMux
    port map (
            O => \N__44907\,
            I => \N__44591\
        );

    \I__10582\ : ClkMux
    port map (
            O => \N__44906\,
            I => \N__44591\
        );

    \I__10581\ : ClkMux
    port map (
            O => \N__44905\,
            I => \N__44591\
        );

    \I__10580\ : ClkMux
    port map (
            O => \N__44904\,
            I => \N__44591\
        );

    \I__10579\ : ClkMux
    port map (
            O => \N__44903\,
            I => \N__44591\
        );

    \I__10578\ : ClkMux
    port map (
            O => \N__44902\,
            I => \N__44591\
        );

    \I__10577\ : ClkMux
    port map (
            O => \N__44901\,
            I => \N__44591\
        );

    \I__10576\ : ClkMux
    port map (
            O => \N__44900\,
            I => \N__44591\
        );

    \I__10575\ : ClkMux
    port map (
            O => \N__44899\,
            I => \N__44591\
        );

    \I__10574\ : ClkMux
    port map (
            O => \N__44898\,
            I => \N__44591\
        );

    \I__10573\ : ClkMux
    port map (
            O => \N__44897\,
            I => \N__44591\
        );

    \I__10572\ : ClkMux
    port map (
            O => \N__44896\,
            I => \N__44591\
        );

    \I__10571\ : ClkMux
    port map (
            O => \N__44895\,
            I => \N__44591\
        );

    \I__10570\ : ClkMux
    port map (
            O => \N__44894\,
            I => \N__44591\
        );

    \I__10569\ : ClkMux
    port map (
            O => \N__44893\,
            I => \N__44591\
        );

    \I__10568\ : ClkMux
    port map (
            O => \N__44892\,
            I => \N__44591\
        );

    \I__10567\ : ClkMux
    port map (
            O => \N__44891\,
            I => \N__44591\
        );

    \I__10566\ : ClkMux
    port map (
            O => \N__44890\,
            I => \N__44591\
        );

    \I__10565\ : ClkMux
    port map (
            O => \N__44889\,
            I => \N__44591\
        );

    \I__10564\ : ClkMux
    port map (
            O => \N__44888\,
            I => \N__44591\
        );

    \I__10563\ : ClkMux
    port map (
            O => \N__44887\,
            I => \N__44591\
        );

    \I__10562\ : ClkMux
    port map (
            O => \N__44886\,
            I => \N__44591\
        );

    \I__10561\ : ClkMux
    port map (
            O => \N__44885\,
            I => \N__44591\
        );

    \I__10560\ : ClkMux
    port map (
            O => \N__44884\,
            I => \N__44591\
        );

    \I__10559\ : ClkMux
    port map (
            O => \N__44883\,
            I => \N__44591\
        );

    \I__10558\ : ClkMux
    port map (
            O => \N__44882\,
            I => \N__44591\
        );

    \I__10557\ : ClkMux
    port map (
            O => \N__44881\,
            I => \N__44591\
        );

    \I__10556\ : ClkMux
    port map (
            O => \N__44880\,
            I => \N__44591\
        );

    \I__10555\ : ClkMux
    port map (
            O => \N__44879\,
            I => \N__44591\
        );

    \I__10554\ : ClkMux
    port map (
            O => \N__44878\,
            I => \N__44591\
        );

    \I__10553\ : ClkMux
    port map (
            O => \N__44877\,
            I => \N__44591\
        );

    \I__10552\ : ClkMux
    port map (
            O => \N__44876\,
            I => \N__44591\
        );

    \I__10551\ : ClkMux
    port map (
            O => \N__44875\,
            I => \N__44591\
        );

    \I__10550\ : ClkMux
    port map (
            O => \N__44874\,
            I => \N__44591\
        );

    \I__10549\ : ClkMux
    port map (
            O => \N__44873\,
            I => \N__44591\
        );

    \I__10548\ : ClkMux
    port map (
            O => \N__44872\,
            I => \N__44591\
        );

    \I__10547\ : ClkMux
    port map (
            O => \N__44871\,
            I => \N__44591\
        );

    \I__10546\ : ClkMux
    port map (
            O => \N__44870\,
            I => \N__44591\
        );

    \I__10545\ : ClkMux
    port map (
            O => \N__44869\,
            I => \N__44591\
        );

    \I__10544\ : ClkMux
    port map (
            O => \N__44868\,
            I => \N__44591\
        );

    \I__10543\ : ClkMux
    port map (
            O => \N__44867\,
            I => \N__44591\
        );

    \I__10542\ : ClkMux
    port map (
            O => \N__44866\,
            I => \N__44591\
        );

    \I__10541\ : ClkMux
    port map (
            O => \N__44865\,
            I => \N__44591\
        );

    \I__10540\ : ClkMux
    port map (
            O => \N__44864\,
            I => \N__44591\
        );

    \I__10539\ : ClkMux
    port map (
            O => \N__44863\,
            I => \N__44591\
        );

    \I__10538\ : ClkMux
    port map (
            O => \N__44862\,
            I => \N__44591\
        );

    \I__10537\ : ClkMux
    port map (
            O => \N__44861\,
            I => \N__44591\
        );

    \I__10536\ : ClkMux
    port map (
            O => \N__44860\,
            I => \N__44591\
        );

    \I__10535\ : ClkMux
    port map (
            O => \N__44859\,
            I => \N__44591\
        );

    \I__10534\ : ClkMux
    port map (
            O => \N__44858\,
            I => \N__44591\
        );

    \I__10533\ : ClkMux
    port map (
            O => \N__44857\,
            I => \N__44591\
        );

    \I__10532\ : ClkMux
    port map (
            O => \N__44856\,
            I => \N__44591\
        );

    \I__10531\ : ClkMux
    port map (
            O => \N__44855\,
            I => \N__44591\
        );

    \I__10530\ : ClkMux
    port map (
            O => \N__44854\,
            I => \N__44591\
        );

    \I__10529\ : ClkMux
    port map (
            O => \N__44853\,
            I => \N__44591\
        );

    \I__10528\ : ClkMux
    port map (
            O => \N__44852\,
            I => \N__44591\
        );

    \I__10527\ : ClkMux
    port map (
            O => \N__44851\,
            I => \N__44591\
        );

    \I__10526\ : ClkMux
    port map (
            O => \N__44850\,
            I => \N__44591\
        );

    \I__10525\ : ClkMux
    port map (
            O => \N__44849\,
            I => \N__44591\
        );

    \I__10524\ : ClkMux
    port map (
            O => \N__44848\,
            I => \N__44591\
        );

    \I__10523\ : ClkMux
    port map (
            O => \N__44847\,
            I => \N__44591\
        );

    \I__10522\ : ClkMux
    port map (
            O => \N__44846\,
            I => \N__44591\
        );

    \I__10521\ : ClkMux
    port map (
            O => \N__44845\,
            I => \N__44591\
        );

    \I__10520\ : ClkMux
    port map (
            O => \N__44844\,
            I => \N__44591\
        );

    \I__10519\ : ClkMux
    port map (
            O => \N__44843\,
            I => \N__44591\
        );

    \I__10518\ : ClkMux
    port map (
            O => \N__44842\,
            I => \N__44591\
        );

    \I__10517\ : ClkMux
    port map (
            O => \N__44841\,
            I => \N__44591\
        );

    \I__10516\ : ClkMux
    port map (
            O => \N__44840\,
            I => \N__44591\
        );

    \I__10515\ : ClkMux
    port map (
            O => \N__44839\,
            I => \N__44591\
        );

    \I__10514\ : ClkMux
    port map (
            O => \N__44838\,
            I => \N__44591\
        );

    \I__10513\ : ClkMux
    port map (
            O => \N__44837\,
            I => \N__44591\
        );

    \I__10512\ : ClkMux
    port map (
            O => \N__44836\,
            I => \N__44591\
        );

    \I__10511\ : ClkMux
    port map (
            O => \N__44835\,
            I => \N__44591\
        );

    \I__10510\ : ClkMux
    port map (
            O => \N__44834\,
            I => \N__44591\
        );

    \I__10509\ : ClkMux
    port map (
            O => \N__44833\,
            I => \N__44591\
        );

    \I__10508\ : ClkMux
    port map (
            O => \N__44832\,
            I => \N__44591\
        );

    \I__10507\ : GlobalMux
    port map (
            O => \N__44591\,
            I => clk_100mhz_0
        );

    \I__10506\ : SRMux
    port map (
            O => \N__44588\,
            I => \N__44584\
        );

    \I__10505\ : SRMux
    port map (
            O => \N__44587\,
            I => \N__44581\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__44584\,
            I => \N__44578\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__44581\,
            I => \N__44573\
        );

    \I__10502\ : Span4Mux_v
    port map (
            O => \N__44578\,
            I => \N__44570\
        );

    \I__10501\ : SRMux
    port map (
            O => \N__44577\,
            I => \N__44567\
        );

    \I__10500\ : SRMux
    port map (
            O => \N__44576\,
            I => \N__44564\
        );

    \I__10499\ : Span4Mux_h
    port map (
            O => \N__44573\,
            I => \N__44561\
        );

    \I__10498\ : Span4Mux_h
    port map (
            O => \N__44570\,
            I => \N__44556\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__44567\,
            I => \N__44556\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__44564\,
            I => \N__44553\
        );

    \I__10495\ : Odrv4
    port map (
            O => \N__44561\,
            I => \phase_controller_inst2.stoper_tr.un1_stoper_state12_1_0_i\
        );

    \I__10494\ : Odrv4
    port map (
            O => \N__44556\,
            I => \phase_controller_inst2.stoper_tr.un1_stoper_state12_1_0_i\
        );

    \I__10493\ : Odrv4
    port map (
            O => \N__44553\,
            I => \phase_controller_inst2.stoper_tr.un1_stoper_state12_1_0_i\
        );

    \I__10492\ : InMux
    port map (
            O => \N__44546\,
            I => \N__44542\
        );

    \I__10491\ : InMux
    port map (
            O => \N__44545\,
            I => \N__44539\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__44542\,
            I => \N__44536\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__44539\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10488\ : Odrv4
    port map (
            O => \N__44536\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10487\ : InMux
    port map (
            O => \N__44531\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__10486\ : InMux
    port map (
            O => \N__44528\,
            I => \N__44524\
        );

    \I__10485\ : InMux
    port map (
            O => \N__44527\,
            I => \N__44521\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__44524\,
            I => \N__44518\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__44521\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__10482\ : Odrv4
    port map (
            O => \N__44518\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__10481\ : InMux
    port map (
            O => \N__44513\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__10480\ : InMux
    port map (
            O => \N__44510\,
            I => \N__44506\
        );

    \I__10479\ : InMux
    port map (
            O => \N__44509\,
            I => \N__44503\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__44506\,
            I => \N__44500\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__44503\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__10476\ : Odrv12
    port map (
            O => \N__44500\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__10475\ : InMux
    port map (
            O => \N__44495\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__10474\ : InMux
    port map (
            O => \N__44492\,
            I => \N__44488\
        );

    \I__10473\ : InMux
    port map (
            O => \N__44491\,
            I => \N__44485\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__44488\,
            I => \N__44482\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__44485\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10470\ : Odrv12
    port map (
            O => \N__44482\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10469\ : InMux
    port map (
            O => \N__44477\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__10468\ : InMux
    port map (
            O => \N__44474\,
            I => \N__44470\
        );

    \I__10467\ : InMux
    port map (
            O => \N__44473\,
            I => \N__44467\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__44470\,
            I => \N__44464\
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__44467\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__10464\ : Odrv4
    port map (
            O => \N__44464\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__10463\ : InMux
    port map (
            O => \N__44459\,
            I => \bfn_18_20_0_\
        );

    \I__10462\ : InMux
    port map (
            O => \N__44456\,
            I => \N__44452\
        );

    \I__10461\ : InMux
    port map (
            O => \N__44455\,
            I => \N__44449\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__44452\,
            I => \N__44446\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__44449\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__10458\ : Odrv4
    port map (
            O => \N__44446\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__10457\ : InMux
    port map (
            O => \N__44441\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__10456\ : InMux
    port map (
            O => \N__44438\,
            I => \N__44434\
        );

    \I__10455\ : InMux
    port map (
            O => \N__44437\,
            I => \N__44431\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__44434\,
            I => \N__44428\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__44431\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10452\ : Odrv4
    port map (
            O => \N__44428\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10451\ : InMux
    port map (
            O => \N__44423\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__10450\ : InMux
    port map (
            O => \N__44420\,
            I => \N__44416\
        );

    \I__10449\ : InMux
    port map (
            O => \N__44419\,
            I => \N__44413\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__44416\,
            I => \N__44410\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__44413\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__10446\ : Odrv4
    port map (
            O => \N__44410\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__10445\ : InMux
    port map (
            O => \N__44405\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__10444\ : InMux
    port map (
            O => \N__44402\,
            I => \N__44398\
        );

    \I__10443\ : InMux
    port map (
            O => \N__44401\,
            I => \N__44395\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__44398\,
            I => \N__44392\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__44395\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__10440\ : Odrv4
    port map (
            O => \N__44392\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__10439\ : InMux
    port map (
            O => \N__44387\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__10438\ : InMux
    port map (
            O => \N__44384\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__10437\ : InMux
    port map (
            O => \N__44381\,
            I => \N__44371\
        );

    \I__10436\ : InMux
    port map (
            O => \N__44380\,
            I => \N__44371\
        );

    \I__10435\ : InMux
    port map (
            O => \N__44379\,
            I => \N__44371\
        );

    \I__10434\ : InMux
    port map (
            O => \N__44378\,
            I => \N__44368\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__44371\,
            I => \N__44364\
        );

    \I__10432\ : LocalMux
    port map (
            O => \N__44368\,
            I => \N__44361\
        );

    \I__10431\ : CascadeMux
    port map (
            O => \N__44367\,
            I => \N__44358\
        );

    \I__10430\ : Span4Mux_h
    port map (
            O => \N__44364\,
            I => \N__44354\
        );

    \I__10429\ : Span4Mux_v
    port map (
            O => \N__44361\,
            I => \N__44351\
        );

    \I__10428\ : InMux
    port map (
            O => \N__44358\,
            I => \N__44346\
        );

    \I__10427\ : InMux
    port map (
            O => \N__44357\,
            I => \N__44346\
        );

    \I__10426\ : Odrv4
    port map (
            O => \N__44354\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10425\ : Odrv4
    port map (
            O => \N__44351\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__44346\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10423\ : CascadeMux
    port map (
            O => \N__44339\,
            I => \N__44328\
        );

    \I__10422\ : CascadeMux
    port map (
            O => \N__44338\,
            I => \N__44323\
        );

    \I__10421\ : InMux
    port map (
            O => \N__44337\,
            I => \N__44308\
        );

    \I__10420\ : InMux
    port map (
            O => \N__44336\,
            I => \N__44305\
        );

    \I__10419\ : InMux
    port map (
            O => \N__44335\,
            I => \N__44302\
        );

    \I__10418\ : InMux
    port map (
            O => \N__44334\,
            I => \N__44299\
        );

    \I__10417\ : InMux
    port map (
            O => \N__44333\,
            I => \N__44296\
        );

    \I__10416\ : InMux
    port map (
            O => \N__44332\,
            I => \N__44293\
        );

    \I__10415\ : InMux
    port map (
            O => \N__44331\,
            I => \N__44290\
        );

    \I__10414\ : InMux
    port map (
            O => \N__44328\,
            I => \N__44285\
        );

    \I__10413\ : InMux
    port map (
            O => \N__44327\,
            I => \N__44285\
        );

    \I__10412\ : InMux
    port map (
            O => \N__44326\,
            I => \N__44282\
        );

    \I__10411\ : InMux
    port map (
            O => \N__44323\,
            I => \N__44275\
        );

    \I__10410\ : InMux
    port map (
            O => \N__44322\,
            I => \N__44275\
        );

    \I__10409\ : InMux
    port map (
            O => \N__44321\,
            I => \N__44275\
        );

    \I__10408\ : InMux
    port map (
            O => \N__44320\,
            I => \N__44272\
        );

    \I__10407\ : InMux
    port map (
            O => \N__44319\,
            I => \N__44267\
        );

    \I__10406\ : InMux
    port map (
            O => \N__44318\,
            I => \N__44267\
        );

    \I__10405\ : InMux
    port map (
            O => \N__44317\,
            I => \N__44262\
        );

    \I__10404\ : InMux
    port map (
            O => \N__44316\,
            I => \N__44262\
        );

    \I__10403\ : InMux
    port map (
            O => \N__44315\,
            I => \N__44259\
        );

    \I__10402\ : InMux
    port map (
            O => \N__44314\,
            I => \N__44254\
        );

    \I__10401\ : InMux
    port map (
            O => \N__44313\,
            I => \N__44254\
        );

    \I__10400\ : InMux
    port map (
            O => \N__44312\,
            I => \N__44249\
        );

    \I__10399\ : InMux
    port map (
            O => \N__44311\,
            I => \N__44249\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__44308\,
            I => \N__44246\
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__44305\,
            I => \N__44243\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__44302\,
            I => \N__44240\
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__44299\,
            I => \N__44235\
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__44296\,
            I => \N__44211\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__44293\,
            I => \N__44205\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__44290\,
            I => \N__44202\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__44285\,
            I => \N__44196\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__44282\,
            I => \N__44193\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__44275\,
            I => \N__44190\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__44272\,
            I => \N__44165\
        );

    \I__10387\ : LocalMux
    port map (
            O => \N__44267\,
            I => \N__44154\
        );

    \I__10386\ : LocalMux
    port map (
            O => \N__44262\,
            I => \N__44147\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__44259\,
            I => \N__44140\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__44254\,
            I => \N__44132\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__44249\,
            I => \N__44126\
        );

    \I__10382\ : Glb2LocalMux
    port map (
            O => \N__44246\,
            I => \N__43874\
        );

    \I__10381\ : Glb2LocalMux
    port map (
            O => \N__44243\,
            I => \N__43874\
        );

    \I__10380\ : Glb2LocalMux
    port map (
            O => \N__44240\,
            I => \N__43874\
        );

    \I__10379\ : SRMux
    port map (
            O => \N__44239\,
            I => \N__43874\
        );

    \I__10378\ : SRMux
    port map (
            O => \N__44238\,
            I => \N__43874\
        );

    \I__10377\ : Glb2LocalMux
    port map (
            O => \N__44235\,
            I => \N__43874\
        );

    \I__10376\ : SRMux
    port map (
            O => \N__44234\,
            I => \N__43874\
        );

    \I__10375\ : SRMux
    port map (
            O => \N__44233\,
            I => \N__43874\
        );

    \I__10374\ : SRMux
    port map (
            O => \N__44232\,
            I => \N__43874\
        );

    \I__10373\ : SRMux
    port map (
            O => \N__44231\,
            I => \N__43874\
        );

    \I__10372\ : SRMux
    port map (
            O => \N__44230\,
            I => \N__43874\
        );

    \I__10371\ : SRMux
    port map (
            O => \N__44229\,
            I => \N__43874\
        );

    \I__10370\ : SRMux
    port map (
            O => \N__44228\,
            I => \N__43874\
        );

    \I__10369\ : SRMux
    port map (
            O => \N__44227\,
            I => \N__43874\
        );

    \I__10368\ : SRMux
    port map (
            O => \N__44226\,
            I => \N__43874\
        );

    \I__10367\ : SRMux
    port map (
            O => \N__44225\,
            I => \N__43874\
        );

    \I__10366\ : SRMux
    port map (
            O => \N__44224\,
            I => \N__43874\
        );

    \I__10365\ : SRMux
    port map (
            O => \N__44223\,
            I => \N__43874\
        );

    \I__10364\ : SRMux
    port map (
            O => \N__44222\,
            I => \N__43874\
        );

    \I__10363\ : SRMux
    port map (
            O => \N__44221\,
            I => \N__43874\
        );

    \I__10362\ : SRMux
    port map (
            O => \N__44220\,
            I => \N__43874\
        );

    \I__10361\ : SRMux
    port map (
            O => \N__44219\,
            I => \N__43874\
        );

    \I__10360\ : SRMux
    port map (
            O => \N__44218\,
            I => \N__43874\
        );

    \I__10359\ : SRMux
    port map (
            O => \N__44217\,
            I => \N__43874\
        );

    \I__10358\ : SRMux
    port map (
            O => \N__44216\,
            I => \N__43874\
        );

    \I__10357\ : SRMux
    port map (
            O => \N__44215\,
            I => \N__43874\
        );

    \I__10356\ : SRMux
    port map (
            O => \N__44214\,
            I => \N__43874\
        );

    \I__10355\ : Glb2LocalMux
    port map (
            O => \N__44211\,
            I => \N__43874\
        );

    \I__10354\ : SRMux
    port map (
            O => \N__44210\,
            I => \N__43874\
        );

    \I__10353\ : SRMux
    port map (
            O => \N__44209\,
            I => \N__43874\
        );

    \I__10352\ : SRMux
    port map (
            O => \N__44208\,
            I => \N__43874\
        );

    \I__10351\ : Glb2LocalMux
    port map (
            O => \N__44205\,
            I => \N__43874\
        );

    \I__10350\ : Glb2LocalMux
    port map (
            O => \N__44202\,
            I => \N__43874\
        );

    \I__10349\ : SRMux
    port map (
            O => \N__44201\,
            I => \N__43874\
        );

    \I__10348\ : SRMux
    port map (
            O => \N__44200\,
            I => \N__43874\
        );

    \I__10347\ : SRMux
    port map (
            O => \N__44199\,
            I => \N__43874\
        );

    \I__10346\ : Glb2LocalMux
    port map (
            O => \N__44196\,
            I => \N__43874\
        );

    \I__10345\ : Glb2LocalMux
    port map (
            O => \N__44193\,
            I => \N__43874\
        );

    \I__10344\ : Glb2LocalMux
    port map (
            O => \N__44190\,
            I => \N__43874\
        );

    \I__10343\ : SRMux
    port map (
            O => \N__44189\,
            I => \N__43874\
        );

    \I__10342\ : SRMux
    port map (
            O => \N__44188\,
            I => \N__43874\
        );

    \I__10341\ : SRMux
    port map (
            O => \N__44187\,
            I => \N__43874\
        );

    \I__10340\ : SRMux
    port map (
            O => \N__44186\,
            I => \N__43874\
        );

    \I__10339\ : SRMux
    port map (
            O => \N__44185\,
            I => \N__43874\
        );

    \I__10338\ : SRMux
    port map (
            O => \N__44184\,
            I => \N__43874\
        );

    \I__10337\ : SRMux
    port map (
            O => \N__44183\,
            I => \N__43874\
        );

    \I__10336\ : SRMux
    port map (
            O => \N__44182\,
            I => \N__43874\
        );

    \I__10335\ : SRMux
    port map (
            O => \N__44181\,
            I => \N__43874\
        );

    \I__10334\ : SRMux
    port map (
            O => \N__44180\,
            I => \N__43874\
        );

    \I__10333\ : SRMux
    port map (
            O => \N__44179\,
            I => \N__43874\
        );

    \I__10332\ : SRMux
    port map (
            O => \N__44178\,
            I => \N__43874\
        );

    \I__10331\ : SRMux
    port map (
            O => \N__44177\,
            I => \N__43874\
        );

    \I__10330\ : SRMux
    port map (
            O => \N__44176\,
            I => \N__43874\
        );

    \I__10329\ : SRMux
    port map (
            O => \N__44175\,
            I => \N__43874\
        );

    \I__10328\ : SRMux
    port map (
            O => \N__44174\,
            I => \N__43874\
        );

    \I__10327\ : SRMux
    port map (
            O => \N__44173\,
            I => \N__43874\
        );

    \I__10326\ : SRMux
    port map (
            O => \N__44172\,
            I => \N__43874\
        );

    \I__10325\ : SRMux
    port map (
            O => \N__44171\,
            I => \N__43874\
        );

    \I__10324\ : SRMux
    port map (
            O => \N__44170\,
            I => \N__43874\
        );

    \I__10323\ : SRMux
    port map (
            O => \N__44169\,
            I => \N__43874\
        );

    \I__10322\ : SRMux
    port map (
            O => \N__44168\,
            I => \N__43874\
        );

    \I__10321\ : Glb2LocalMux
    port map (
            O => \N__44165\,
            I => \N__43874\
        );

    \I__10320\ : SRMux
    port map (
            O => \N__44164\,
            I => \N__43874\
        );

    \I__10319\ : SRMux
    port map (
            O => \N__44163\,
            I => \N__43874\
        );

    \I__10318\ : SRMux
    port map (
            O => \N__44162\,
            I => \N__43874\
        );

    \I__10317\ : SRMux
    port map (
            O => \N__44161\,
            I => \N__43874\
        );

    \I__10316\ : SRMux
    port map (
            O => \N__44160\,
            I => \N__43874\
        );

    \I__10315\ : SRMux
    port map (
            O => \N__44159\,
            I => \N__43874\
        );

    \I__10314\ : SRMux
    port map (
            O => \N__44158\,
            I => \N__43874\
        );

    \I__10313\ : SRMux
    port map (
            O => \N__44157\,
            I => \N__43874\
        );

    \I__10312\ : Glb2LocalMux
    port map (
            O => \N__44154\,
            I => \N__43874\
        );

    \I__10311\ : SRMux
    port map (
            O => \N__44153\,
            I => \N__43874\
        );

    \I__10310\ : SRMux
    port map (
            O => \N__44152\,
            I => \N__43874\
        );

    \I__10309\ : SRMux
    port map (
            O => \N__44151\,
            I => \N__43874\
        );

    \I__10308\ : SRMux
    port map (
            O => \N__44150\,
            I => \N__43874\
        );

    \I__10307\ : Glb2LocalMux
    port map (
            O => \N__44147\,
            I => \N__43874\
        );

    \I__10306\ : SRMux
    port map (
            O => \N__44146\,
            I => \N__43874\
        );

    \I__10305\ : SRMux
    port map (
            O => \N__44145\,
            I => \N__43874\
        );

    \I__10304\ : SRMux
    port map (
            O => \N__44144\,
            I => \N__43874\
        );

    \I__10303\ : SRMux
    port map (
            O => \N__44143\,
            I => \N__43874\
        );

    \I__10302\ : Glb2LocalMux
    port map (
            O => \N__44140\,
            I => \N__43874\
        );

    \I__10301\ : SRMux
    port map (
            O => \N__44139\,
            I => \N__43874\
        );

    \I__10300\ : SRMux
    port map (
            O => \N__44138\,
            I => \N__43874\
        );

    \I__10299\ : SRMux
    port map (
            O => \N__44137\,
            I => \N__43874\
        );

    \I__10298\ : SRMux
    port map (
            O => \N__44136\,
            I => \N__43874\
        );

    \I__10297\ : SRMux
    port map (
            O => \N__44135\,
            I => \N__43874\
        );

    \I__10296\ : Glb2LocalMux
    port map (
            O => \N__44132\,
            I => \N__43874\
        );

    \I__10295\ : SRMux
    port map (
            O => \N__44131\,
            I => \N__43874\
        );

    \I__10294\ : SRMux
    port map (
            O => \N__44130\,
            I => \N__43874\
        );

    \I__10293\ : SRMux
    port map (
            O => \N__44129\,
            I => \N__43874\
        );

    \I__10292\ : Glb2LocalMux
    port map (
            O => \N__44126\,
            I => \N__43874\
        );

    \I__10291\ : SRMux
    port map (
            O => \N__44125\,
            I => \N__43874\
        );

    \I__10290\ : SRMux
    port map (
            O => \N__44124\,
            I => \N__43874\
        );

    \I__10289\ : SRMux
    port map (
            O => \N__44123\,
            I => \N__43874\
        );

    \I__10288\ : SRMux
    port map (
            O => \N__44122\,
            I => \N__43874\
        );

    \I__10287\ : SRMux
    port map (
            O => \N__44121\,
            I => \N__43874\
        );

    \I__10286\ : SRMux
    port map (
            O => \N__44120\,
            I => \N__43874\
        );

    \I__10285\ : SRMux
    port map (
            O => \N__44119\,
            I => \N__43874\
        );

    \I__10284\ : SRMux
    port map (
            O => \N__44118\,
            I => \N__43874\
        );

    \I__10283\ : SRMux
    port map (
            O => \N__44117\,
            I => \N__43874\
        );

    \I__10282\ : SRMux
    port map (
            O => \N__44116\,
            I => \N__43874\
        );

    \I__10281\ : SRMux
    port map (
            O => \N__44115\,
            I => \N__43874\
        );

    \I__10280\ : SRMux
    port map (
            O => \N__44114\,
            I => \N__43874\
        );

    \I__10279\ : SRMux
    port map (
            O => \N__44113\,
            I => \N__43874\
        );

    \I__10278\ : SRMux
    port map (
            O => \N__44112\,
            I => \N__43874\
        );

    \I__10277\ : SRMux
    port map (
            O => \N__44111\,
            I => \N__43874\
        );

    \I__10276\ : SRMux
    port map (
            O => \N__44110\,
            I => \N__43874\
        );

    \I__10275\ : SRMux
    port map (
            O => \N__44109\,
            I => \N__43874\
        );

    \I__10274\ : SRMux
    port map (
            O => \N__44108\,
            I => \N__43874\
        );

    \I__10273\ : SRMux
    port map (
            O => \N__44107\,
            I => \N__43874\
        );

    \I__10272\ : SRMux
    port map (
            O => \N__44106\,
            I => \N__43874\
        );

    \I__10271\ : SRMux
    port map (
            O => \N__44105\,
            I => \N__43874\
        );

    \I__10270\ : SRMux
    port map (
            O => \N__44104\,
            I => \N__43874\
        );

    \I__10269\ : SRMux
    port map (
            O => \N__44103\,
            I => \N__43874\
        );

    \I__10268\ : GlobalMux
    port map (
            O => \N__43874\,
            I => \N__43871\
        );

    \I__10267\ : gio2CtrlBuf
    port map (
            O => \N__43871\,
            I => red_c_g
        );

    \I__10266\ : InMux
    port map (
            O => \N__43868\,
            I => \N__43865\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__43865\,
            I => \N__43861\
        );

    \I__10264\ : CascadeMux
    port map (
            O => \N__43864\,
            I => \N__43857\
        );

    \I__10263\ : Span4Mux_h
    port map (
            O => \N__43861\,
            I => \N__43852\
        );

    \I__10262\ : InMux
    port map (
            O => \N__43860\,
            I => \N__43843\
        );

    \I__10261\ : InMux
    port map (
            O => \N__43857\,
            I => \N__43843\
        );

    \I__10260\ : InMux
    port map (
            O => \N__43856\,
            I => \N__43843\
        );

    \I__10259\ : InMux
    port map (
            O => \N__43855\,
            I => \N__43843\
        );

    \I__10258\ : Odrv4
    port map (
            O => \N__43852\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__43843\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__10256\ : InMux
    port map (
            O => \N__43838\,
            I => \N__43834\
        );

    \I__10255\ : CascadeMux
    port map (
            O => \N__43837\,
            I => \N__43829\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__43834\,
            I => \N__43823\
        );

    \I__10253\ : CascadeMux
    port map (
            O => \N__43833\,
            I => \N__43820\
        );

    \I__10252\ : CascadeMux
    port map (
            O => \N__43832\,
            I => \N__43816\
        );

    \I__10251\ : InMux
    port map (
            O => \N__43829\,
            I => \N__43809\
        );

    \I__10250\ : InMux
    port map (
            O => \N__43828\,
            I => \N__43809\
        );

    \I__10249\ : InMux
    port map (
            O => \N__43827\,
            I => \N__43809\
        );

    \I__10248\ : InMux
    port map (
            O => \N__43826\,
            I => \N__43806\
        );

    \I__10247\ : Span4Mux_v
    port map (
            O => \N__43823\,
            I => \N__43803\
        );

    \I__10246\ : InMux
    port map (
            O => \N__43820\,
            I => \N__43796\
        );

    \I__10245\ : InMux
    port map (
            O => \N__43819\,
            I => \N__43796\
        );

    \I__10244\ : InMux
    port map (
            O => \N__43816\,
            I => \N__43796\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__43809\,
            I => \N__43793\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__43806\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10241\ : Odrv4
    port map (
            O => \N__43803\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__43796\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10239\ : Odrv4
    port map (
            O => \N__43793\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10238\ : InMux
    port map (
            O => \N__43784\,
            I => \N__43781\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__43781\,
            I => \N__43774\
        );

    \I__10236\ : InMux
    port map (
            O => \N__43780\,
            I => \N__43765\
        );

    \I__10235\ : InMux
    port map (
            O => \N__43779\,
            I => \N__43765\
        );

    \I__10234\ : InMux
    port map (
            O => \N__43778\,
            I => \N__43765\
        );

    \I__10233\ : InMux
    port map (
            O => \N__43777\,
            I => \N__43765\
        );

    \I__10232\ : Span4Mux_v
    port map (
            O => \N__43774\,
            I => \N__43760\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__43765\,
            I => \N__43760\
        );

    \I__10230\ : Span4Mux_h
    port map (
            O => \N__43760\,
            I => \N__43756\
        );

    \I__10229\ : InMux
    port map (
            O => \N__43759\,
            I => \N__43753\
        );

    \I__10228\ : Span4Mux_h
    port map (
            O => \N__43756\,
            I => \N__43750\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__43753\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__10226\ : Odrv4
    port map (
            O => \N__43750\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__10225\ : CEMux
    port map (
            O => \N__43745\,
            I => \N__43740\
        );

    \I__10224\ : CEMux
    port map (
            O => \N__43744\,
            I => \N__43737\
        );

    \I__10223\ : CEMux
    port map (
            O => \N__43743\,
            I => \N__43732\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__43740\,
            I => \N__43729\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__43737\,
            I => \N__43726\
        );

    \I__10220\ : CEMux
    port map (
            O => \N__43736\,
            I => \N__43723\
        );

    \I__10219\ : CEMux
    port map (
            O => \N__43735\,
            I => \N__43720\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__43732\,
            I => \N__43717\
        );

    \I__10217\ : Span4Mux_v
    port map (
            O => \N__43729\,
            I => \N__43714\
        );

    \I__10216\ : Span4Mux_v
    port map (
            O => \N__43726\,
            I => \N__43711\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__43723\,
            I => \N__43708\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__43720\,
            I => \N__43705\
        );

    \I__10213\ : Span4Mux_h
    port map (
            O => \N__43717\,
            I => \N__43702\
        );

    \I__10212\ : Span4Mux_v
    port map (
            O => \N__43714\,
            I => \N__43699\
        );

    \I__10211\ : Span4Mux_v
    port map (
            O => \N__43711\,
            I => \N__43694\
        );

    \I__10210\ : Span4Mux_h
    port map (
            O => \N__43708\,
            I => \N__43694\
        );

    \I__10209\ : Span4Mux_v
    port map (
            O => \N__43705\,
            I => \N__43691\
        );

    \I__10208\ : Odrv4
    port map (
            O => \N__43702\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0\
        );

    \I__10207\ : Odrv4
    port map (
            O => \N__43699\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0\
        );

    \I__10206\ : Odrv4
    port map (
            O => \N__43694\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0\
        );

    \I__10205\ : Odrv4
    port map (
            O => \N__43691\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0\
        );

    \I__10204\ : InMux
    port map (
            O => \N__43682\,
            I => \N__43678\
        );

    \I__10203\ : InMux
    port map (
            O => \N__43681\,
            I => \N__43675\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__43678\,
            I => \N__43672\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__43675\,
            I => \N__43668\
        );

    \I__10200\ : Span4Mux_v
    port map (
            O => \N__43672\,
            I => \N__43665\
        );

    \I__10199\ : InMux
    port map (
            O => \N__43671\,
            I => \N__43662\
        );

    \I__10198\ : Span4Mux_h
    port map (
            O => \N__43668\,
            I => \N__43659\
        );

    \I__10197\ : Span4Mux_h
    port map (
            O => \N__43665\,
            I => \N__43656\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__43662\,
            I => \N__43651\
        );

    \I__10195\ : Span4Mux_v
    port map (
            O => \N__43659\,
            I => \N__43651\
        );

    \I__10194\ : Odrv4
    port map (
            O => \N__43656\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10193\ : Odrv4
    port map (
            O => \N__43651\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10192\ : CascadeMux
    port map (
            O => \N__43646\,
            I => \N__43643\
        );

    \I__10191\ : InMux
    port map (
            O => \N__43643\,
            I => \N__43640\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__43640\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__10189\ : InMux
    port map (
            O => \N__43637\,
            I => \N__43633\
        );

    \I__10188\ : InMux
    port map (
            O => \N__43636\,
            I => \N__43630\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__43633\,
            I => \N__43627\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__43630\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__10185\ : Odrv4
    port map (
            O => \N__43627\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__10184\ : InMux
    port map (
            O => \N__43622\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__10183\ : CascadeMux
    port map (
            O => \N__43619\,
            I => \N__43616\
        );

    \I__10182\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43613\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__43613\,
            I => \N__43610\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__43610\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84ADZ0\
        );

    \I__10179\ : InMux
    port map (
            O => \N__43607\,
            I => \N__43603\
        );

    \I__10178\ : InMux
    port map (
            O => \N__43606\,
            I => \N__43600\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__43603\,
            I => \N__43597\
        );

    \I__10176\ : LocalMux
    port map (
            O => \N__43600\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__10175\ : Odrv4
    port map (
            O => \N__43597\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__10174\ : InMux
    port map (
            O => \N__43592\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__10173\ : InMux
    port map (
            O => \N__43589\,
            I => \N__43585\
        );

    \I__10172\ : InMux
    port map (
            O => \N__43588\,
            I => \N__43582\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__43585\,
            I => \N__43579\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__43582\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__10169\ : Odrv4
    port map (
            O => \N__43579\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__10168\ : InMux
    port map (
            O => \N__43574\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__10167\ : InMux
    port map (
            O => \N__43571\,
            I => \N__43568\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__43568\,
            I => \N__43565\
        );

    \I__10165\ : Span4Mux_v
    port map (
            O => \N__43565\,
            I => \N__43562\
        );

    \I__10164\ : Odrv4
    port map (
            O => \N__43562\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__10163\ : CascadeMux
    port map (
            O => \N__43559\,
            I => \N__43556\
        );

    \I__10162\ : InMux
    port map (
            O => \N__43556\,
            I => \N__43553\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__43553\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__10160\ : InMux
    port map (
            O => \N__43550\,
            I => \N__43547\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__43547\,
            I => \N__43544\
        );

    \I__10158\ : Span4Mux_v
    port map (
            O => \N__43544\,
            I => \N__43541\
        );

    \I__10157\ : Odrv4
    port map (
            O => \N__43541\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__10156\ : CascadeMux
    port map (
            O => \N__43538\,
            I => \N__43535\
        );

    \I__10155\ : InMux
    port map (
            O => \N__43535\,
            I => \N__43532\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__43532\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__10153\ : InMux
    port map (
            O => \N__43529\,
            I => \N__43526\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__43526\,
            I => \N__43523\
        );

    \I__10151\ : Odrv12
    port map (
            O => \N__43523\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__10150\ : CascadeMux
    port map (
            O => \N__43520\,
            I => \N__43517\
        );

    \I__10149\ : InMux
    port map (
            O => \N__43517\,
            I => \N__43514\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__43514\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__10147\ : InMux
    port map (
            O => \N__43511\,
            I => \N__43508\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__43508\,
            I => \N__43505\
        );

    \I__10145\ : Span4Mux_v
    port map (
            O => \N__43505\,
            I => \N__43502\
        );

    \I__10144\ : Odrv4
    port map (
            O => \N__43502\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__10143\ : CascadeMux
    port map (
            O => \N__43499\,
            I => \N__43496\
        );

    \I__10142\ : InMux
    port map (
            O => \N__43496\,
            I => \N__43493\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__43493\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__10140\ : CascadeMux
    port map (
            O => \N__43490\,
            I => \N__43487\
        );

    \I__10139\ : InMux
    port map (
            O => \N__43487\,
            I => \N__43484\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__43484\,
            I => \N__43481\
        );

    \I__10137\ : Span4Mux_h
    port map (
            O => \N__43481\,
            I => \N__43478\
        );

    \I__10136\ : Odrv4
    port map (
            O => \N__43478\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__10135\ : InMux
    port map (
            O => \N__43475\,
            I => \N__43472\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__43472\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\
        );

    \I__10133\ : InMux
    port map (
            O => \N__43469\,
            I => \N__43466\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__43466\,
            I => \N__43463\
        );

    \I__10131\ : Span4Mux_h
    port map (
            O => \N__43463\,
            I => \N__43460\
        );

    \I__10130\ : Odrv4
    port map (
            O => \N__43460\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__10129\ : CascadeMux
    port map (
            O => \N__43457\,
            I => \N__43454\
        );

    \I__10128\ : InMux
    port map (
            O => \N__43454\,
            I => \N__43451\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__43451\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\
        );

    \I__10126\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43445\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__43445\,
            I => \N__43442\
        );

    \I__10124\ : Odrv12
    port map (
            O => \N__43442\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__10123\ : CascadeMux
    port map (
            O => \N__43439\,
            I => \N__43436\
        );

    \I__10122\ : InMux
    port map (
            O => \N__43436\,
            I => \N__43433\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__43433\,
            I => \N__43430\
        );

    \I__10120\ : Odrv4
    port map (
            O => \N__43430\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\
        );

    \I__10119\ : InMux
    port map (
            O => \N__43427\,
            I => \N__43424\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__43424\,
            I => \N__43421\
        );

    \I__10117\ : Span4Mux_v
    port map (
            O => \N__43421\,
            I => \N__43418\
        );

    \I__10116\ : Odrv4
    port map (
            O => \N__43418\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__10115\ : CascadeMux
    port map (
            O => \N__43415\,
            I => \N__43412\
        );

    \I__10114\ : InMux
    port map (
            O => \N__43412\,
            I => \N__43409\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__43409\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\
        );

    \I__10112\ : CascadeMux
    port map (
            O => \N__43406\,
            I => \N__43403\
        );

    \I__10111\ : InMux
    port map (
            O => \N__43403\,
            I => \N__43400\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__43400\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__10109\ : CascadeMux
    port map (
            O => \N__43397\,
            I => \N__43394\
        );

    \I__10108\ : InMux
    port map (
            O => \N__43394\,
            I => \N__43391\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__43391\,
            I => \N__43388\
        );

    \I__10106\ : Odrv4
    port map (
            O => \N__43388\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__10105\ : InMux
    port map (
            O => \N__43385\,
            I => \N__43382\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__43382\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__10103\ : InMux
    port map (
            O => \N__43379\,
            I => \N__43376\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__43376\,
            I => \N__43373\
        );

    \I__10101\ : Span4Mux_h
    port map (
            O => \N__43373\,
            I => \N__43370\
        );

    \I__10100\ : Odrv4
    port map (
            O => \N__43370\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__10099\ : CascadeMux
    port map (
            O => \N__43367\,
            I => \N__43364\
        );

    \I__10098\ : InMux
    port map (
            O => \N__43364\,
            I => \N__43361\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__43361\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__10096\ : InMux
    port map (
            O => \N__43358\,
            I => \N__43355\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__43355\,
            I => \N__43352\
        );

    \I__10094\ : Span4Mux_h
    port map (
            O => \N__43352\,
            I => \N__43349\
        );

    \I__10093\ : Odrv4
    port map (
            O => \N__43349\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__10092\ : CascadeMux
    port map (
            O => \N__43346\,
            I => \N__43343\
        );

    \I__10091\ : InMux
    port map (
            O => \N__43343\,
            I => \N__43340\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__43340\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__10089\ : InMux
    port map (
            O => \N__43337\,
            I => \N__43334\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__43334\,
            I => \N__43331\
        );

    \I__10087\ : Span4Mux_v
    port map (
            O => \N__43331\,
            I => \N__43328\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__43328\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__10085\ : CascadeMux
    port map (
            O => \N__43325\,
            I => \N__43322\
        );

    \I__10084\ : InMux
    port map (
            O => \N__43322\,
            I => \N__43319\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__43319\,
            I => \N__43316\
        );

    \I__10082\ : Odrv4
    port map (
            O => \N__43316\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__10081\ : InMux
    port map (
            O => \N__43313\,
            I => \N__43310\
        );

    \I__10080\ : LocalMux
    port map (
            O => \N__43310\,
            I => \N__43307\
        );

    \I__10079\ : Span4Mux_h
    port map (
            O => \N__43307\,
            I => \N__43304\
        );

    \I__10078\ : Span4Mux_h
    port map (
            O => \N__43304\,
            I => \N__43301\
        );

    \I__10077\ : Odrv4
    port map (
            O => \N__43301\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__10076\ : CascadeMux
    port map (
            O => \N__43298\,
            I => \N__43295\
        );

    \I__10075\ : InMux
    port map (
            O => \N__43295\,
            I => \N__43292\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__43292\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__10073\ : InMux
    port map (
            O => \N__43289\,
            I => \N__43286\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__43286\,
            I => \N__43283\
        );

    \I__10071\ : Odrv12
    port map (
            O => \N__43283\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__10070\ : CascadeMux
    port map (
            O => \N__43280\,
            I => \N__43277\
        );

    \I__10069\ : InMux
    port map (
            O => \N__43277\,
            I => \N__43274\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__43274\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__10067\ : CascadeMux
    port map (
            O => \N__43271\,
            I => \N__43268\
        );

    \I__10066\ : InMux
    port map (
            O => \N__43268\,
            I => \N__43265\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__43265\,
            I => \N__43262\
        );

    \I__10064\ : Odrv12
    port map (
            O => \N__43262\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__10063\ : InMux
    port map (
            O => \N__43259\,
            I => \N__43256\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__43256\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__10061\ : InMux
    port map (
            O => \N__43253\,
            I => \N__43249\
        );

    \I__10060\ : InMux
    port map (
            O => \N__43252\,
            I => \N__43246\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__43249\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__43246\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10057\ : InMux
    port map (
            O => \N__43241\,
            I => \N__43238\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__43238\,
            I => \N__43235\
        );

    \I__10055\ : Odrv4
    port map (
            O => \N__43235\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__10054\ : CascadeMux
    port map (
            O => \N__43232\,
            I => \N__43229\
        );

    \I__10053\ : InMux
    port map (
            O => \N__43229\,
            I => \N__43226\
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__43226\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__10051\ : InMux
    port map (
            O => \N__43223\,
            I => \N__43220\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__43220\,
            I => \N__43217\
        );

    \I__10049\ : Odrv4
    port map (
            O => \N__43217\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__10048\ : InMux
    port map (
            O => \N__43214\,
            I => \N__43210\
        );

    \I__10047\ : InMux
    port map (
            O => \N__43213\,
            I => \N__43207\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__43210\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__43207\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10044\ : CascadeMux
    port map (
            O => \N__43202\,
            I => \N__43199\
        );

    \I__10043\ : InMux
    port map (
            O => \N__43199\,
            I => \N__43196\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__43196\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__10041\ : InMux
    port map (
            O => \N__43193\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__10040\ : InMux
    port map (
            O => \N__43190\,
            I => \N__43185\
        );

    \I__10039\ : InMux
    port map (
            O => \N__43189\,
            I => \N__43182\
        );

    \I__10038\ : CascadeMux
    port map (
            O => \N__43188\,
            I => \N__43175\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__43185\,
            I => \N__43171\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__43182\,
            I => \N__43168\
        );

    \I__10035\ : InMux
    port map (
            O => \N__43181\,
            I => \N__43155\
        );

    \I__10034\ : InMux
    port map (
            O => \N__43180\,
            I => \N__43155\
        );

    \I__10033\ : InMux
    port map (
            O => \N__43179\,
            I => \N__43155\
        );

    \I__10032\ : InMux
    port map (
            O => \N__43178\,
            I => \N__43155\
        );

    \I__10031\ : InMux
    port map (
            O => \N__43175\,
            I => \N__43155\
        );

    \I__10030\ : InMux
    port map (
            O => \N__43174\,
            I => \N__43155\
        );

    \I__10029\ : Odrv4
    port map (
            O => \N__43171\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10028\ : Odrv12
    port map (
            O => \N__43168\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__43155\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10026\ : InMux
    port map (
            O => \N__43148\,
            I => \N__43145\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__43145\,
            I => \N__43140\
        );

    \I__10024\ : CascadeMux
    port map (
            O => \N__43144\,
            I => \N__43136\
        );

    \I__10023\ : CascadeMux
    port map (
            O => \N__43143\,
            I => \N__43133\
        );

    \I__10022\ : Span4Mux_v
    port map (
            O => \N__43140\,
            I => \N__43128\
        );

    \I__10021\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43119\
        );

    \I__10020\ : InMux
    port map (
            O => \N__43136\,
            I => \N__43119\
        );

    \I__10019\ : InMux
    port map (
            O => \N__43133\,
            I => \N__43119\
        );

    \I__10018\ : InMux
    port map (
            O => \N__43132\,
            I => \N__43119\
        );

    \I__10017\ : InMux
    port map (
            O => \N__43131\,
            I => \N__43116\
        );

    \I__10016\ : Sp12to4
    port map (
            O => \N__43128\,
            I => \N__43111\
        );

    \I__10015\ : LocalMux
    port map (
            O => \N__43119\,
            I => \N__43111\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__43116\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10013\ : Odrv12
    port map (
            O => \N__43111\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10012\ : InMux
    port map (
            O => \N__43106\,
            I => \N__43103\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__43103\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0\
        );

    \I__10010\ : CascadeMux
    port map (
            O => \N__43100\,
            I => \N__43097\
        );

    \I__10009\ : InMux
    port map (
            O => \N__43097\,
            I => \N__43094\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__43094\,
            I => \N__43091\
        );

    \I__10007\ : Span4Mux_v
    port map (
            O => \N__43091\,
            I => \N__43088\
        );

    \I__10006\ : Odrv4
    port map (
            O => \N__43088\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__10005\ : InMux
    port map (
            O => \N__43085\,
            I => \N__43082\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__43082\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__10003\ : InMux
    port map (
            O => \N__43079\,
            I => \N__43076\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__43076\,
            I => \N__43073\
        );

    \I__10001\ : Odrv4
    port map (
            O => \N__43073\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__10000\ : CascadeMux
    port map (
            O => \N__43070\,
            I => \N__43067\
        );

    \I__9999\ : InMux
    port map (
            O => \N__43067\,
            I => \N__43064\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__43064\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__9997\ : InMux
    port map (
            O => \N__43061\,
            I => \N__43058\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__43058\,
            I => \N__43055\
        );

    \I__9995\ : Span4Mux_v
    port map (
            O => \N__43055\,
            I => \N__43052\
        );

    \I__9994\ : Odrv4
    port map (
            O => \N__43052\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__9993\ : CascadeMux
    port map (
            O => \N__43049\,
            I => \N__43046\
        );

    \I__9992\ : InMux
    port map (
            O => \N__43046\,
            I => \N__43043\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__43043\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__9990\ : InMux
    port map (
            O => \N__43040\,
            I => \N__43037\
        );

    \I__9989\ : LocalMux
    port map (
            O => \N__43037\,
            I => \N__43034\
        );

    \I__9988\ : Odrv12
    port map (
            O => \N__43034\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__9987\ : InMux
    port map (
            O => \N__43031\,
            I => \N__43027\
        );

    \I__9986\ : InMux
    port map (
            O => \N__43030\,
            I => \N__43024\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__43027\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__43024\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__9983\ : InMux
    port map (
            O => \N__43019\,
            I => \N__43016\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__43016\,
            I => \N__43013\
        );

    \I__9981\ : Odrv4
    port map (
            O => \N__43013\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__9980\ : CascadeMux
    port map (
            O => \N__43010\,
            I => \N__43007\
        );

    \I__9979\ : InMux
    port map (
            O => \N__43007\,
            I => \N__43004\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__43004\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__9977\ : InMux
    port map (
            O => \N__43001\,
            I => \N__42998\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__42998\,
            I => \N__42995\
        );

    \I__9975\ : Odrv4
    port map (
            O => \N__42995\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__9974\ : InMux
    port map (
            O => \N__42992\,
            I => \N__42988\
        );

    \I__9973\ : InMux
    port map (
            O => \N__42991\,
            I => \N__42985\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__42988\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__42985\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__9970\ : CascadeMux
    port map (
            O => \N__42980\,
            I => \N__42977\
        );

    \I__9969\ : InMux
    port map (
            O => \N__42977\,
            I => \N__42974\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__42974\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__9967\ : InMux
    port map (
            O => \N__42971\,
            I => \N__42968\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__42968\,
            I => \N__42965\
        );

    \I__9965\ : Span4Mux_v
    port map (
            O => \N__42965\,
            I => \N__42962\
        );

    \I__9964\ : Odrv4
    port map (
            O => \N__42962\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__9963\ : InMux
    port map (
            O => \N__42959\,
            I => \N__42955\
        );

    \I__9962\ : InMux
    port map (
            O => \N__42958\,
            I => \N__42952\
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__42955\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__42952\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__42947\,
            I => \N__42944\
        );

    \I__9958\ : InMux
    port map (
            O => \N__42944\,
            I => \N__42941\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__42941\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__9956\ : CascadeMux
    port map (
            O => \N__42938\,
            I => \N__42935\
        );

    \I__9955\ : InMux
    port map (
            O => \N__42935\,
            I => \N__42932\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__42932\,
            I => \N__42929\
        );

    \I__9953\ : Odrv4
    port map (
            O => \N__42929\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__9952\ : InMux
    port map (
            O => \N__42926\,
            I => \N__42922\
        );

    \I__9951\ : InMux
    port map (
            O => \N__42925\,
            I => \N__42919\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__42922\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__42919\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__9948\ : InMux
    port map (
            O => \N__42914\,
            I => \N__42911\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__42911\,
            I => \N__42908\
        );

    \I__9946\ : Odrv4
    port map (
            O => \N__42908\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__9945\ : InMux
    port map (
            O => \N__42905\,
            I => \N__42902\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__42902\,
            I => \N__42899\
        );

    \I__9943\ : Odrv4
    port map (
            O => \N__42899\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__9942\ : InMux
    port map (
            O => \N__42896\,
            I => \N__42892\
        );

    \I__9941\ : InMux
    port map (
            O => \N__42895\,
            I => \N__42889\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__42892\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__42889\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__9938\ : CascadeMux
    port map (
            O => \N__42884\,
            I => \N__42881\
        );

    \I__9937\ : InMux
    port map (
            O => \N__42881\,
            I => \N__42878\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__42878\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__9935\ : CascadeMux
    port map (
            O => \N__42875\,
            I => \N__42872\
        );

    \I__9934\ : InMux
    port map (
            O => \N__42872\,
            I => \N__42869\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__42869\,
            I => \N__42866\
        );

    \I__9932\ : Span4Mux_h
    port map (
            O => \N__42866\,
            I => \N__42863\
        );

    \I__9931\ : Odrv4
    port map (
            O => \N__42863\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__9930\ : InMux
    port map (
            O => \N__42860\,
            I => \N__42856\
        );

    \I__9929\ : InMux
    port map (
            O => \N__42859\,
            I => \N__42853\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__42856\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__42853\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__9926\ : InMux
    port map (
            O => \N__42848\,
            I => \N__42845\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__42845\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__9924\ : InMux
    port map (
            O => \N__42842\,
            I => \N__42838\
        );

    \I__9923\ : InMux
    port map (
            O => \N__42841\,
            I => \N__42835\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__42838\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__42835\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9920\ : InMux
    port map (
            O => \N__42830\,
            I => \N__42827\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__42827\,
            I => \N__42824\
        );

    \I__9918\ : Odrv4
    port map (
            O => \N__42824\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__9917\ : CascadeMux
    port map (
            O => \N__42821\,
            I => \N__42818\
        );

    \I__9916\ : InMux
    port map (
            O => \N__42818\,
            I => \N__42815\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__42815\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__9914\ : CascadeMux
    port map (
            O => \N__42812\,
            I => \N__42809\
        );

    \I__9913\ : InMux
    port map (
            O => \N__42809\,
            I => \N__42806\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__42806\,
            I => \N__42803\
        );

    \I__9911\ : Odrv12
    port map (
            O => \N__42803\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__9910\ : InMux
    port map (
            O => \N__42800\,
            I => \N__42796\
        );

    \I__9909\ : InMux
    port map (
            O => \N__42799\,
            I => \N__42793\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__42796\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__42793\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9906\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42785\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__42785\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__9904\ : CascadeMux
    port map (
            O => \N__42782\,
            I => \N__42779\
        );

    \I__9903\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42776\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__42776\,
            I => \N__42773\
        );

    \I__9901\ : Span4Mux_h
    port map (
            O => \N__42773\,
            I => \N__42770\
        );

    \I__9900\ : Span4Mux_v
    port map (
            O => \N__42770\,
            I => \N__42767\
        );

    \I__9899\ : Odrv4
    port map (
            O => \N__42767\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__9898\ : CascadeMux
    port map (
            O => \N__42764\,
            I => \N__42761\
        );

    \I__9897\ : InMux
    port map (
            O => \N__42761\,
            I => \N__42757\
        );

    \I__9896\ : InMux
    port map (
            O => \N__42760\,
            I => \N__42754\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__42757\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__42754\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__9893\ : InMux
    port map (
            O => \N__42749\,
            I => \N__42746\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__42746\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__9891\ : InMux
    port map (
            O => \N__42743\,
            I => \N__42740\
        );

    \I__9890\ : LocalMux
    port map (
            O => \N__42740\,
            I => \N__42737\
        );

    \I__9889\ : Span4Mux_h
    port map (
            O => \N__42737\,
            I => \N__42734\
        );

    \I__9888\ : Span4Mux_v
    port map (
            O => \N__42734\,
            I => \N__42731\
        );

    \I__9887\ : Odrv4
    port map (
            O => \N__42731\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__9886\ : InMux
    port map (
            O => \N__42728\,
            I => \N__42724\
        );

    \I__9885\ : InMux
    port map (
            O => \N__42727\,
            I => \N__42721\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__42724\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__42721\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__9882\ : CascadeMux
    port map (
            O => \N__42716\,
            I => \N__42713\
        );

    \I__9881\ : InMux
    port map (
            O => \N__42713\,
            I => \N__42710\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__42710\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__9879\ : InMux
    port map (
            O => \N__42707\,
            I => \N__42704\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__42704\,
            I => \N__42701\
        );

    \I__9877\ : Span4Mux_v
    port map (
            O => \N__42701\,
            I => \N__42698\
        );

    \I__9876\ : Odrv4
    port map (
            O => \N__42698\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__9875\ : InMux
    port map (
            O => \N__42695\,
            I => \N__42691\
        );

    \I__9874\ : InMux
    port map (
            O => \N__42694\,
            I => \N__42688\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__42691\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__42688\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__9871\ : CascadeMux
    port map (
            O => \N__42683\,
            I => \N__42680\
        );

    \I__9870\ : InMux
    port map (
            O => \N__42680\,
            I => \N__42677\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__42677\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__9868\ : InMux
    port map (
            O => \N__42674\,
            I => \N__42671\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__42671\,
            I => \N__42668\
        );

    \I__9866\ : Span4Mux_h
    port map (
            O => \N__42668\,
            I => \N__42665\
        );

    \I__9865\ : Odrv4
    port map (
            O => \N__42665\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__9864\ : InMux
    port map (
            O => \N__42662\,
            I => \N__42658\
        );

    \I__9863\ : InMux
    port map (
            O => \N__42661\,
            I => \N__42655\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__42658\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__42655\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__9860\ : CascadeMux
    port map (
            O => \N__42650\,
            I => \N__42647\
        );

    \I__9859\ : InMux
    port map (
            O => \N__42647\,
            I => \N__42644\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__42644\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__9857\ : InMux
    port map (
            O => \N__42641\,
            I => \N__42638\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__42638\,
            I => \N__42635\
        );

    \I__9855\ : Span4Mux_v
    port map (
            O => \N__42635\,
            I => \N__42632\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__42632\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__9853\ : InMux
    port map (
            O => \N__42629\,
            I => \N__42625\
        );

    \I__9852\ : InMux
    port map (
            O => \N__42628\,
            I => \N__42622\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__42625\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__42622\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__9849\ : CascadeMux
    port map (
            O => \N__42617\,
            I => \N__42614\
        );

    \I__9848\ : InMux
    port map (
            O => \N__42614\,
            I => \N__42611\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__42611\,
            I => \N__42608\
        );

    \I__9846\ : Odrv4
    port map (
            O => \N__42608\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__9845\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42601\
        );

    \I__9844\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42598\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__42601\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__42598\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__9841\ : InMux
    port map (
            O => \N__42593\,
            I => \N__42590\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__42590\,
            I => \N__42587\
        );

    \I__9839\ : Span4Mux_h
    port map (
            O => \N__42587\,
            I => \N__42584\
        );

    \I__9838\ : Odrv4
    port map (
            O => \N__42584\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__9837\ : CascadeMux
    port map (
            O => \N__42581\,
            I => \N__42578\
        );

    \I__9836\ : InMux
    port map (
            O => \N__42578\,
            I => \N__42575\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__42575\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__9834\ : InMux
    port map (
            O => \N__42572\,
            I => \N__42569\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__42569\,
            I => \N__42566\
        );

    \I__9832\ : Span4Mux_v
    port map (
            O => \N__42566\,
            I => \N__42563\
        );

    \I__9831\ : Odrv4
    port map (
            O => \N__42563\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__9830\ : InMux
    port map (
            O => \N__42560\,
            I => \N__42556\
        );

    \I__9829\ : InMux
    port map (
            O => \N__42559\,
            I => \N__42553\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__42556\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__42553\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__9826\ : CascadeMux
    port map (
            O => \N__42548\,
            I => \N__42545\
        );

    \I__9825\ : InMux
    port map (
            O => \N__42545\,
            I => \N__42542\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__42542\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__9823\ : CascadeMux
    port map (
            O => \N__42539\,
            I => \N__42536\
        );

    \I__9822\ : InMux
    port map (
            O => \N__42536\,
            I => \N__42531\
        );

    \I__9821\ : CascadeMux
    port map (
            O => \N__42535\,
            I => \N__42528\
        );

    \I__9820\ : InMux
    port map (
            O => \N__42534\,
            I => \N__42525\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__42531\,
            I => \N__42522\
        );

    \I__9818\ : InMux
    port map (
            O => \N__42528\,
            I => \N__42518\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__42525\,
            I => \N__42515\
        );

    \I__9816\ : Span4Mux_h
    port map (
            O => \N__42522\,
            I => \N__42512\
        );

    \I__9815\ : InMux
    port map (
            O => \N__42521\,
            I => \N__42509\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__42518\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__9813\ : Odrv12
    port map (
            O => \N__42515\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__9812\ : Odrv4
    port map (
            O => \N__42512\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__42509\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__9810\ : InMux
    port map (
            O => \N__42500\,
            I => \N__42495\
        );

    \I__9809\ : InMux
    port map (
            O => \N__42499\,
            I => \N__42489\
        );

    \I__9808\ : InMux
    port map (
            O => \N__42498\,
            I => \N__42489\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__42495\,
            I => \N__42485\
        );

    \I__9806\ : InMux
    port map (
            O => \N__42494\,
            I => \N__42482\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__42489\,
            I => \N__42479\
        );

    \I__9804\ : InMux
    port map (
            O => \N__42488\,
            I => \N__42476\
        );

    \I__9803\ : Span4Mux_v
    port map (
            O => \N__42485\,
            I => \N__42473\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__42482\,
            I => \N__42470\
        );

    \I__9801\ : Span4Mux_h
    port map (
            O => \N__42479\,
            I => \N__42467\
        );

    \I__9800\ : LocalMux
    port map (
            O => \N__42476\,
            I => \elapsed_time_ns_1_RNIFG4DM1_0_16\
        );

    \I__9799\ : Odrv4
    port map (
            O => \N__42473\,
            I => \elapsed_time_ns_1_RNIFG4DM1_0_16\
        );

    \I__9798\ : Odrv12
    port map (
            O => \N__42470\,
            I => \elapsed_time_ns_1_RNIFG4DM1_0_16\
        );

    \I__9797\ : Odrv4
    port map (
            O => \N__42467\,
            I => \elapsed_time_ns_1_RNIFG4DM1_0_16\
        );

    \I__9796\ : InMux
    port map (
            O => \N__42458\,
            I => \N__42441\
        );

    \I__9795\ : InMux
    port map (
            O => \N__42457\,
            I => \N__42441\
        );

    \I__9794\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42441\
        );

    \I__9793\ : InMux
    port map (
            O => \N__42455\,
            I => \N__42441\
        );

    \I__9792\ : InMux
    port map (
            O => \N__42454\,
            I => \N__42430\
        );

    \I__9791\ : InMux
    port map (
            O => \N__42453\,
            I => \N__42430\
        );

    \I__9790\ : InMux
    port map (
            O => \N__42452\,
            I => \N__42430\
        );

    \I__9789\ : InMux
    port map (
            O => \N__42451\,
            I => \N__42430\
        );

    \I__9788\ : InMux
    port map (
            O => \N__42450\,
            I => \N__42430\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__42441\,
            I => \N__42424\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__42430\,
            I => \N__42424\
        );

    \I__9785\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42421\
        );

    \I__9784\ : Span4Mux_v
    port map (
            O => \N__42424\,
            I => \N__42418\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__42421\,
            I => \phase_controller_inst1.stoper_tr.N_241\
        );

    \I__9782\ : Odrv4
    port map (
            O => \N__42418\,
            I => \phase_controller_inst1.stoper_tr.N_241\
        );

    \I__9781\ : CascadeMux
    port map (
            O => \N__42413\,
            I => \N__42409\
        );

    \I__9780\ : InMux
    port map (
            O => \N__42412\,
            I => \N__42406\
        );

    \I__9779\ : InMux
    port map (
            O => \N__42409\,
            I => \N__42403\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__42406\,
            I => \N__42400\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__42403\,
            I => \N__42397\
        );

    \I__9776\ : Span4Mux_h
    port map (
            O => \N__42400\,
            I => \N__42393\
        );

    \I__9775\ : Span4Mux_v
    port map (
            O => \N__42397\,
            I => \N__42390\
        );

    \I__9774\ : InMux
    port map (
            O => \N__42396\,
            I => \N__42387\
        );

    \I__9773\ : Odrv4
    port map (
            O => \N__42393\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__9772\ : Odrv4
    port map (
            O => \N__42390\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__42387\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__9770\ : InMux
    port map (
            O => \N__42380\,
            I => \N__42376\
        );

    \I__9769\ : InMux
    port map (
            O => \N__42379\,
            I => \N__42373\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__42376\,
            I => \N__42366\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__42373\,
            I => \N__42366\
        );

    \I__9766\ : CascadeMux
    port map (
            O => \N__42372\,
            I => \N__42362\
        );

    \I__9765\ : InMux
    port map (
            O => \N__42371\,
            I => \N__42359\
        );

    \I__9764\ : Span4Mux_v
    port map (
            O => \N__42366\,
            I => \N__42356\
        );

    \I__9763\ : InMux
    port map (
            O => \N__42365\,
            I => \N__42351\
        );

    \I__9762\ : InMux
    port map (
            O => \N__42362\,
            I => \N__42351\
        );

    \I__9761\ : LocalMux
    port map (
            O => \N__42359\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19\
        );

    \I__9760\ : Odrv4
    port map (
            O => \N__42356\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__42351\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19\
        );

    \I__9758\ : InMux
    port map (
            O => \N__42344\,
            I => \N__42340\
        );

    \I__9757\ : InMux
    port map (
            O => \N__42343\,
            I => \N__42337\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__42340\,
            I => \N__42334\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__42337\,
            I => \N__42331\
        );

    \I__9754\ : Span4Mux_h
    port map (
            O => \N__42334\,
            I => \N__42325\
        );

    \I__9753\ : Span4Mux_v
    port map (
            O => \N__42331\,
            I => \N__42325\
        );

    \I__9752\ : InMux
    port map (
            O => \N__42330\,
            I => \N__42320\
        );

    \I__9751\ : Span4Mux_h
    port map (
            O => \N__42325\,
            I => \N__42317\
        );

    \I__9750\ : InMux
    port map (
            O => \N__42324\,
            I => \N__42312\
        );

    \I__9749\ : InMux
    port map (
            O => \N__42323\,
            I => \N__42312\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__42320\,
            I => \elapsed_time_ns_1_RNIHI4DM1_0_18\
        );

    \I__9747\ : Odrv4
    port map (
            O => \N__42317\,
            I => \elapsed_time_ns_1_RNIHI4DM1_0_18\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__42312\,
            I => \elapsed_time_ns_1_RNIHI4DM1_0_18\
        );

    \I__9745\ : InMux
    port map (
            O => \N__42305\,
            I => \N__42300\
        );

    \I__9744\ : InMux
    port map (
            O => \N__42304\,
            I => \N__42297\
        );

    \I__9743\ : InMux
    port map (
            O => \N__42303\,
            I => \N__42294\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__42300\,
            I => \N__42291\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__42297\,
            I => \N__42286\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__42294\,
            I => \N__42281\
        );

    \I__9739\ : Span4Mux_h
    port map (
            O => \N__42291\,
            I => \N__42281\
        );

    \I__9738\ : InMux
    port map (
            O => \N__42290\,
            I => \N__42276\
        );

    \I__9737\ : InMux
    port map (
            O => \N__42289\,
            I => \N__42276\
        );

    \I__9736\ : Odrv4
    port map (
            O => \N__42286\,
            I => \elapsed_time_ns_1_RNIGH4DM1_0_17\
        );

    \I__9735\ : Odrv4
    port map (
            O => \N__42281\,
            I => \elapsed_time_ns_1_RNIGH4DM1_0_17\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__42276\,
            I => \elapsed_time_ns_1_RNIGH4DM1_0_17\
        );

    \I__9733\ : CascadeMux
    port map (
            O => \N__42269\,
            I => \N__42261\
        );

    \I__9732\ : CascadeMux
    port map (
            O => \N__42268\,
            I => \N__42257\
        );

    \I__9731\ : CascadeMux
    port map (
            O => \N__42267\,
            I => \N__42253\
        );

    \I__9730\ : InMux
    port map (
            O => \N__42266\,
            I => \N__42233\
        );

    \I__9729\ : InMux
    port map (
            O => \N__42265\,
            I => \N__42233\
        );

    \I__9728\ : InMux
    port map (
            O => \N__42264\,
            I => \N__42233\
        );

    \I__9727\ : InMux
    port map (
            O => \N__42261\,
            I => \N__42233\
        );

    \I__9726\ : InMux
    port map (
            O => \N__42260\,
            I => \N__42233\
        );

    \I__9725\ : InMux
    port map (
            O => \N__42257\,
            I => \N__42228\
        );

    \I__9724\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42228\
        );

    \I__9723\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42222\
        );

    \I__9722\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42222\
        );

    \I__9721\ : InMux
    port map (
            O => \N__42251\,
            I => \N__42215\
        );

    \I__9720\ : InMux
    port map (
            O => \N__42250\,
            I => \N__42215\
        );

    \I__9719\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42215\
        );

    \I__9718\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42204\
        );

    \I__9717\ : InMux
    port map (
            O => \N__42247\,
            I => \N__42204\
        );

    \I__9716\ : InMux
    port map (
            O => \N__42246\,
            I => \N__42204\
        );

    \I__9715\ : InMux
    port map (
            O => \N__42245\,
            I => \N__42204\
        );

    \I__9714\ : InMux
    port map (
            O => \N__42244\,
            I => \N__42204\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__42233\,
            I => \N__42199\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__42228\,
            I => \N__42199\
        );

    \I__9711\ : CascadeMux
    port map (
            O => \N__42227\,
            I => \N__42191\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__42222\,
            I => \N__42176\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__42215\,
            I => \N__42171\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__42204\,
            I => \N__42171\
        );

    \I__9707\ : Span4Mux_h
    port map (
            O => \N__42199\,
            I => \N__42168\
        );

    \I__9706\ : InMux
    port map (
            O => \N__42198\,
            I => \N__42158\
        );

    \I__9705\ : InMux
    port map (
            O => \N__42197\,
            I => \N__42158\
        );

    \I__9704\ : InMux
    port map (
            O => \N__42196\,
            I => \N__42158\
        );

    \I__9703\ : InMux
    port map (
            O => \N__42195\,
            I => \N__42141\
        );

    \I__9702\ : InMux
    port map (
            O => \N__42194\,
            I => \N__42141\
        );

    \I__9701\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42141\
        );

    \I__9700\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42141\
        );

    \I__9699\ : InMux
    port map (
            O => \N__42189\,
            I => \N__42141\
        );

    \I__9698\ : InMux
    port map (
            O => \N__42188\,
            I => \N__42141\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42187\,
            I => \N__42141\
        );

    \I__9696\ : InMux
    port map (
            O => \N__42186\,
            I => \N__42141\
        );

    \I__9695\ : InMux
    port map (
            O => \N__42185\,
            I => \N__42126\
        );

    \I__9694\ : InMux
    port map (
            O => \N__42184\,
            I => \N__42126\
        );

    \I__9693\ : InMux
    port map (
            O => \N__42183\,
            I => \N__42126\
        );

    \I__9692\ : InMux
    port map (
            O => \N__42182\,
            I => \N__42126\
        );

    \I__9691\ : InMux
    port map (
            O => \N__42181\,
            I => \N__42126\
        );

    \I__9690\ : InMux
    port map (
            O => \N__42180\,
            I => \N__42126\
        );

    \I__9689\ : InMux
    port map (
            O => \N__42179\,
            I => \N__42126\
        );

    \I__9688\ : Span4Mux_v
    port map (
            O => \N__42176\,
            I => \N__42123\
        );

    \I__9687\ : Span4Mux_h
    port map (
            O => \N__42171\,
            I => \N__42120\
        );

    \I__9686\ : Span4Mux_v
    port map (
            O => \N__42168\,
            I => \N__42117\
        );

    \I__9685\ : InMux
    port map (
            O => \N__42167\,
            I => \N__42114\
        );

    \I__9684\ : InMux
    port map (
            O => \N__42166\,
            I => \N__42109\
        );

    \I__9683\ : InMux
    port map (
            O => \N__42165\,
            I => \N__42109\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__42158\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__42141\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__42126\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9679\ : Odrv4
    port map (
            O => \N__42123\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9678\ : Odrv4
    port map (
            O => \N__42120\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9677\ : Odrv4
    port map (
            O => \N__42117\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__42114\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__42109\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9674\ : CascadeMux
    port map (
            O => \N__42092\,
            I => \N__42082\
        );

    \I__9673\ : CascadeMux
    port map (
            O => \N__42091\,
            I => \N__42079\
        );

    \I__9672\ : CascadeMux
    port map (
            O => \N__42090\,
            I => \N__42076\
        );

    \I__9671\ : CascadeMux
    port map (
            O => \N__42089\,
            I => \N__42063\
        );

    \I__9670\ : InMux
    port map (
            O => \N__42088\,
            I => \N__42043\
        );

    \I__9669\ : InMux
    port map (
            O => \N__42087\,
            I => \N__42043\
        );

    \I__9668\ : InMux
    port map (
            O => \N__42086\,
            I => \N__42043\
        );

    \I__9667\ : InMux
    port map (
            O => \N__42085\,
            I => \N__42043\
        );

    \I__9666\ : InMux
    port map (
            O => \N__42082\,
            I => \N__42043\
        );

    \I__9665\ : InMux
    port map (
            O => \N__42079\,
            I => \N__42043\
        );

    \I__9664\ : InMux
    port map (
            O => \N__42076\,
            I => \N__42043\
        );

    \I__9663\ : InMux
    port map (
            O => \N__42075\,
            I => \N__42043\
        );

    \I__9662\ : CascadeMux
    port map (
            O => \N__42074\,
            I => \N__42039\
        );

    \I__9661\ : InMux
    port map (
            O => \N__42073\,
            I => \N__42029\
        );

    \I__9660\ : InMux
    port map (
            O => \N__42072\,
            I => \N__42029\
        );

    \I__9659\ : InMux
    port map (
            O => \N__42071\,
            I => \N__42029\
        );

    \I__9658\ : InMux
    port map (
            O => \N__42070\,
            I => \N__42029\
        );

    \I__9657\ : InMux
    port map (
            O => \N__42069\,
            I => \N__42026\
        );

    \I__9656\ : InMux
    port map (
            O => \N__42068\,
            I => \N__42010\
        );

    \I__9655\ : InMux
    port map (
            O => \N__42067\,
            I => \N__42010\
        );

    \I__9654\ : InMux
    port map (
            O => \N__42066\,
            I => \N__42010\
        );

    \I__9653\ : InMux
    port map (
            O => \N__42063\,
            I => \N__42010\
        );

    \I__9652\ : InMux
    port map (
            O => \N__42062\,
            I => \N__42010\
        );

    \I__9651\ : InMux
    port map (
            O => \N__42061\,
            I => \N__42010\
        );

    \I__9650\ : InMux
    port map (
            O => \N__42060\,
            I => \N__42010\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__42043\,
            I => \N__42003\
        );

    \I__9648\ : InMux
    port map (
            O => \N__42042\,
            I => \N__41996\
        );

    \I__9647\ : InMux
    port map (
            O => \N__42039\,
            I => \N__41996\
        );

    \I__9646\ : InMux
    port map (
            O => \N__42038\,
            I => \N__41996\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__42029\,
            I => \N__41993\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__42026\,
            I => \N__41990\
        );

    \I__9643\ : InMux
    port map (
            O => \N__42025\,
            I => \N__41987\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__42010\,
            I => \N__41984\
        );

    \I__9641\ : InMux
    port map (
            O => \N__42009\,
            I => \N__41981\
        );

    \I__9640\ : InMux
    port map (
            O => \N__42008\,
            I => \N__41978\
        );

    \I__9639\ : InMux
    port map (
            O => \N__42007\,
            I => \N__41973\
        );

    \I__9638\ : InMux
    port map (
            O => \N__42006\,
            I => \N__41973\
        );

    \I__9637\ : Span4Mux_h
    port map (
            O => \N__42003\,
            I => \N__41970\
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__41996\,
            I => \N__41961\
        );

    \I__9635\ : Span4Mux_v
    port map (
            O => \N__41993\,
            I => \N__41961\
        );

    \I__9634\ : Span4Mux_h
    port map (
            O => \N__41990\,
            I => \N__41961\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__41987\,
            I => \N__41961\
        );

    \I__9632\ : Span4Mux_h
    port map (
            O => \N__41984\,
            I => \N__41952\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__41981\,
            I => \N__41952\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__41978\,
            I => \N__41952\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__41973\,
            I => \N__41952\
        );

    \I__9628\ : Odrv4
    port map (
            O => \N__41970\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0Z0Z_15\
        );

    \I__9627\ : Odrv4
    port map (
            O => \N__41961\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0Z0Z_15\
        );

    \I__9626\ : Odrv4
    port map (
            O => \N__41952\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0Z0Z_15\
        );

    \I__9625\ : CEMux
    port map (
            O => \N__41945\,
            I => \N__41942\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__41942\,
            I => \N__41938\
        );

    \I__9623\ : CEMux
    port map (
            O => \N__41941\,
            I => \N__41935\
        );

    \I__9622\ : Span4Mux_v
    port map (
            O => \N__41938\,
            I => \N__41931\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__41935\,
            I => \N__41928\
        );

    \I__9620\ : CEMux
    port map (
            O => \N__41934\,
            I => \N__41925\
        );

    \I__9619\ : Span4Mux_h
    port map (
            O => \N__41931\,
            I => \N__41920\
        );

    \I__9618\ : Span4Mux_v
    port map (
            O => \N__41928\,
            I => \N__41920\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__41925\,
            I => \N__41917\
        );

    \I__9616\ : Span4Mux_v
    port map (
            O => \N__41920\,
            I => \N__41914\
        );

    \I__9615\ : Span4Mux_h
    port map (
            O => \N__41917\,
            I => \N__41911\
        );

    \I__9614\ : Odrv4
    port map (
            O => \N__41914\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa_0\
        );

    \I__9613\ : Odrv4
    port map (
            O => \N__41911\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa_0\
        );

    \I__9612\ : InMux
    port map (
            O => \N__41906\,
            I => \N__41903\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__41903\,
            I => \N__41900\
        );

    \I__9610\ : Span4Mux_h
    port map (
            O => \N__41900\,
            I => \N__41897\
        );

    \I__9609\ : Span4Mux_v
    port map (
            O => \N__41897\,
            I => \N__41894\
        );

    \I__9608\ : Span4Mux_v
    port map (
            O => \N__41894\,
            I => \N__41891\
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__41891\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__9606\ : InMux
    port map (
            O => \N__41888\,
            I => \N__41885\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__41885\,
            I => \N__41882\
        );

    \I__9604\ : Span4Mux_v
    port map (
            O => \N__41882\,
            I => \N__41877\
        );

    \I__9603\ : InMux
    port map (
            O => \N__41881\,
            I => \N__41874\
        );

    \I__9602\ : InMux
    port map (
            O => \N__41880\,
            I => \N__41871\
        );

    \I__9601\ : Sp12to4
    port map (
            O => \N__41877\,
            I => \N__41866\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__41874\,
            I => \N__41866\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__41871\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__9598\ : Odrv12
    port map (
            O => \N__41866\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__9597\ : CascadeMux
    port map (
            O => \N__41861\,
            I => \N__41858\
        );

    \I__9596\ : InMux
    port map (
            O => \N__41858\,
            I => \N__41855\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__41855\,
            I => \N__41852\
        );

    \I__9594\ : Odrv4
    port map (
            O => \N__41852\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__9593\ : InMux
    port map (
            O => \N__41849\,
            I => \N__41845\
        );

    \I__9592\ : InMux
    port map (
            O => \N__41848\,
            I => \N__41842\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__41845\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__41842\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__9589\ : InMux
    port map (
            O => \N__41837\,
            I => \N__41834\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__41834\,
            I => \N__41831\
        );

    \I__9587\ : Span4Mux_h
    port map (
            O => \N__41831\,
            I => \N__41828\
        );

    \I__9586\ : Odrv4
    port map (
            O => \N__41828\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__9585\ : CascadeMux
    port map (
            O => \N__41825\,
            I => \N__41822\
        );

    \I__9584\ : InMux
    port map (
            O => \N__41822\,
            I => \N__41819\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__41819\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__9582\ : InMux
    port map (
            O => \N__41816\,
            I => \N__41778\
        );

    \I__9581\ : InMux
    port map (
            O => \N__41815\,
            I => \N__41778\
        );

    \I__9580\ : InMux
    port map (
            O => \N__41814\,
            I => \N__41778\
        );

    \I__9579\ : InMux
    port map (
            O => \N__41813\,
            I => \N__41778\
        );

    \I__9578\ : InMux
    port map (
            O => \N__41812\,
            I => \N__41769\
        );

    \I__9577\ : InMux
    port map (
            O => \N__41811\,
            I => \N__41769\
        );

    \I__9576\ : InMux
    port map (
            O => \N__41810\,
            I => \N__41769\
        );

    \I__9575\ : InMux
    port map (
            O => \N__41809\,
            I => \N__41769\
        );

    \I__9574\ : InMux
    port map (
            O => \N__41808\,
            I => \N__41764\
        );

    \I__9573\ : InMux
    port map (
            O => \N__41807\,
            I => \N__41764\
        );

    \I__9572\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41755\
        );

    \I__9571\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41755\
        );

    \I__9570\ : InMux
    port map (
            O => \N__41804\,
            I => \N__41755\
        );

    \I__9569\ : InMux
    port map (
            O => \N__41803\,
            I => \N__41755\
        );

    \I__9568\ : InMux
    port map (
            O => \N__41802\,
            I => \N__41746\
        );

    \I__9567\ : InMux
    port map (
            O => \N__41801\,
            I => \N__41746\
        );

    \I__9566\ : InMux
    port map (
            O => \N__41800\,
            I => \N__41746\
        );

    \I__9565\ : InMux
    port map (
            O => \N__41799\,
            I => \N__41746\
        );

    \I__9564\ : InMux
    port map (
            O => \N__41798\,
            I => \N__41737\
        );

    \I__9563\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41737\
        );

    \I__9562\ : InMux
    port map (
            O => \N__41796\,
            I => \N__41737\
        );

    \I__9561\ : InMux
    port map (
            O => \N__41795\,
            I => \N__41737\
        );

    \I__9560\ : InMux
    port map (
            O => \N__41794\,
            I => \N__41728\
        );

    \I__9559\ : InMux
    port map (
            O => \N__41793\,
            I => \N__41728\
        );

    \I__9558\ : InMux
    port map (
            O => \N__41792\,
            I => \N__41728\
        );

    \I__9557\ : InMux
    port map (
            O => \N__41791\,
            I => \N__41728\
        );

    \I__9556\ : InMux
    port map (
            O => \N__41790\,
            I => \N__41719\
        );

    \I__9555\ : InMux
    port map (
            O => \N__41789\,
            I => \N__41719\
        );

    \I__9554\ : InMux
    port map (
            O => \N__41788\,
            I => \N__41719\
        );

    \I__9553\ : InMux
    port map (
            O => \N__41787\,
            I => \N__41719\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__41778\,
            I => \N__41714\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__41769\,
            I => \N__41714\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__41764\,
            I => \N__41711\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__41755\,
            I => \N__41704\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__41746\,
            I => \N__41704\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__41737\,
            I => \N__41704\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__41728\,
            I => \N__41699\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__41719\,
            I => \N__41699\
        );

    \I__9544\ : Span4Mux_h
    port map (
            O => \N__41714\,
            I => \N__41696\
        );

    \I__9543\ : Span4Mux_h
    port map (
            O => \N__41711\,
            I => \N__41693\
        );

    \I__9542\ : Span4Mux_v
    port map (
            O => \N__41704\,
            I => \N__41686\
        );

    \I__9541\ : Span4Mux_v
    port map (
            O => \N__41699\,
            I => \N__41686\
        );

    \I__9540\ : Span4Mux_v
    port map (
            O => \N__41696\,
            I => \N__41686\
        );

    \I__9539\ : Odrv4
    port map (
            O => \N__41693\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9538\ : Odrv4
    port map (
            O => \N__41686\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9537\ : InMux
    port map (
            O => \N__41681\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__9536\ : CascadeMux
    port map (
            O => \N__41678\,
            I => \N__41675\
        );

    \I__9535\ : InMux
    port map (
            O => \N__41675\,
            I => \N__41672\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__41672\,
            I => \N__41668\
        );

    \I__9533\ : InMux
    port map (
            O => \N__41671\,
            I => \N__41665\
        );

    \I__9532\ : Span4Mux_h
    port map (
            O => \N__41668\,
            I => \N__41662\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__41665\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__9530\ : Odrv4
    port map (
            O => \N__41662\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__9529\ : CEMux
    port map (
            O => \N__41657\,
            I => \N__41652\
        );

    \I__9528\ : CEMux
    port map (
            O => \N__41656\,
            I => \N__41649\
        );

    \I__9527\ : CEMux
    port map (
            O => \N__41655\,
            I => \N__41646\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__41652\,
            I => \N__41642\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__41649\,
            I => \N__41639\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__41646\,
            I => \N__41636\
        );

    \I__9523\ : CEMux
    port map (
            O => \N__41645\,
            I => \N__41633\
        );

    \I__9522\ : Span4Mux_v
    port map (
            O => \N__41642\,
            I => \N__41630\
        );

    \I__9521\ : Span4Mux_h
    port map (
            O => \N__41639\,
            I => \N__41627\
        );

    \I__9520\ : Span4Mux_h
    port map (
            O => \N__41636\,
            I => \N__41624\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__41633\,
            I => \N__41621\
        );

    \I__9518\ : Span4Mux_v
    port map (
            O => \N__41630\,
            I => \N__41618\
        );

    \I__9517\ : Span4Mux_v
    port map (
            O => \N__41627\,
            I => \N__41615\
        );

    \I__9516\ : Span4Mux_h
    port map (
            O => \N__41624\,
            I => \N__41612\
        );

    \I__9515\ : Span4Mux_h
    port map (
            O => \N__41621\,
            I => \N__41609\
        );

    \I__9514\ : Odrv4
    port map (
            O => \N__41618\,
            I => \delay_measurement_inst.delay_tr_timer.N_435_i\
        );

    \I__9513\ : Odrv4
    port map (
            O => \N__41615\,
            I => \delay_measurement_inst.delay_tr_timer.N_435_i\
        );

    \I__9512\ : Odrv4
    port map (
            O => \N__41612\,
            I => \delay_measurement_inst.delay_tr_timer.N_435_i\
        );

    \I__9511\ : Odrv4
    port map (
            O => \N__41609\,
            I => \delay_measurement_inst.delay_tr_timer.N_435_i\
        );

    \I__9510\ : CascadeMux
    port map (
            O => \N__41600\,
            I => \N__41597\
        );

    \I__9509\ : InMux
    port map (
            O => \N__41597\,
            I => \N__41593\
        );

    \I__9508\ : InMux
    port map (
            O => \N__41596\,
            I => \N__41589\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__41593\,
            I => \N__41586\
        );

    \I__9506\ : InMux
    port map (
            O => \N__41592\,
            I => \N__41582\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__41589\,
            I => \N__41577\
        );

    \I__9504\ : Span4Mux_h
    port map (
            O => \N__41586\,
            I => \N__41577\
        );

    \I__9503\ : InMux
    port map (
            O => \N__41585\,
            I => \N__41574\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__41582\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__9501\ : Odrv4
    port map (
            O => \N__41577\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__41574\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__9499\ : InMux
    port map (
            O => \N__41567\,
            I => \N__41563\
        );

    \I__9498\ : InMux
    port map (
            O => \N__41566\,
            I => \N__41560\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__41563\,
            I => \N__41557\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__41560\,
            I => \N__41554\
        );

    \I__9495\ : Span4Mux_h
    port map (
            O => \N__41557\,
            I => \N__41548\
        );

    \I__9494\ : Span4Mux_h
    port map (
            O => \N__41554\,
            I => \N__41545\
        );

    \I__9493\ : InMux
    port map (
            O => \N__41553\,
            I => \N__41540\
        );

    \I__9492\ : InMux
    port map (
            O => \N__41552\,
            I => \N__41540\
        );

    \I__9491\ : InMux
    port map (
            O => \N__41551\,
            I => \N__41537\
        );

    \I__9490\ : Odrv4
    port map (
            O => \N__41548\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__9489\ : Odrv4
    port map (
            O => \N__41545\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__41540\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__9487\ : LocalMux
    port map (
            O => \N__41537\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__9486\ : CascadeMux
    port map (
            O => \N__41528\,
            I => \N__41524\
        );

    \I__9485\ : InMux
    port map (
            O => \N__41527\,
            I => \N__41521\
        );

    \I__9484\ : InMux
    port map (
            O => \N__41524\,
            I => \N__41518\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__41521\,
            I => \N__41512\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__41518\,
            I => \N__41512\
        );

    \I__9481\ : InMux
    port map (
            O => \N__41517\,
            I => \N__41508\
        );

    \I__9480\ : Span4Mux_v
    port map (
            O => \N__41512\,
            I => \N__41505\
        );

    \I__9479\ : InMux
    port map (
            O => \N__41511\,
            I => \N__41502\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__41508\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__9477\ : Odrv4
    port map (
            O => \N__41505\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__41502\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__9475\ : CascadeMux
    port map (
            O => \N__41495\,
            I => \N__41492\
        );

    \I__9474\ : InMux
    port map (
            O => \N__41492\,
            I => \N__41488\
        );

    \I__9473\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41484\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__41488\,
            I => \N__41481\
        );

    \I__9471\ : InMux
    port map (
            O => \N__41487\,
            I => \N__41478\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__41484\,
            I => \N__41473\
        );

    \I__9469\ : Span4Mux_h
    port map (
            O => \N__41481\,
            I => \N__41473\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__41478\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__9467\ : Odrv4
    port map (
            O => \N__41473\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__9466\ : InMux
    port map (
            O => \N__41468\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__9465\ : InMux
    port map (
            O => \N__41465\,
            I => \N__41458\
        );

    \I__9464\ : InMux
    port map (
            O => \N__41464\,
            I => \N__41458\
        );

    \I__9463\ : InMux
    port map (
            O => \N__41463\,
            I => \N__41455\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__41458\,
            I => \N__41452\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__41455\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__9460\ : Odrv4
    port map (
            O => \N__41452\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__9459\ : InMux
    port map (
            O => \N__41447\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__9458\ : CascadeMux
    port map (
            O => \N__41444\,
            I => \N__41440\
        );

    \I__9457\ : CascadeMux
    port map (
            O => \N__41443\,
            I => \N__41437\
        );

    \I__9456\ : InMux
    port map (
            O => \N__41440\,
            I => \N__41431\
        );

    \I__9455\ : InMux
    port map (
            O => \N__41437\,
            I => \N__41431\
        );

    \I__9454\ : InMux
    port map (
            O => \N__41436\,
            I => \N__41428\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__41431\,
            I => \N__41425\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__41428\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__41425\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__9450\ : InMux
    port map (
            O => \N__41420\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__9449\ : InMux
    port map (
            O => \N__41417\,
            I => \N__41413\
        );

    \I__9448\ : CascadeMux
    port map (
            O => \N__41416\,
            I => \N__41410\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__41413\,
            I => \N__41406\
        );

    \I__9446\ : InMux
    port map (
            O => \N__41410\,
            I => \N__41403\
        );

    \I__9445\ : InMux
    port map (
            O => \N__41409\,
            I => \N__41400\
        );

    \I__9444\ : Span4Mux_v
    port map (
            O => \N__41406\,
            I => \N__41395\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__41403\,
            I => \N__41395\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__41400\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__9441\ : Odrv4
    port map (
            O => \N__41395\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__9440\ : InMux
    port map (
            O => \N__41390\,
            I => \bfn_18_10_0_\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__41387\,
            I => \N__41384\
        );

    \I__9438\ : InMux
    port map (
            O => \N__41384\,
            I => \N__41380\
        );

    \I__9437\ : InMux
    port map (
            O => \N__41383\,
            I => \N__41376\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__41380\,
            I => \N__41373\
        );

    \I__9435\ : InMux
    port map (
            O => \N__41379\,
            I => \N__41370\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__41376\,
            I => \N__41365\
        );

    \I__9433\ : Span4Mux_v
    port map (
            O => \N__41373\,
            I => \N__41365\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__41370\,
            I => \N__41362\
        );

    \I__9431\ : Odrv4
    port map (
            O => \N__41365\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__9430\ : Odrv4
    port map (
            O => \N__41362\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__9429\ : InMux
    port map (
            O => \N__41357\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__9428\ : CascadeMux
    port map (
            O => \N__41354\,
            I => \N__41350\
        );

    \I__9427\ : CascadeMux
    port map (
            O => \N__41353\,
            I => \N__41347\
        );

    \I__9426\ : InMux
    port map (
            O => \N__41350\,
            I => \N__41341\
        );

    \I__9425\ : InMux
    port map (
            O => \N__41347\,
            I => \N__41341\
        );

    \I__9424\ : InMux
    port map (
            O => \N__41346\,
            I => \N__41338\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__41341\,
            I => \N__41335\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__41338\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__9421\ : Odrv4
    port map (
            O => \N__41335\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__9420\ : InMux
    port map (
            O => \N__41330\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__9419\ : InMux
    port map (
            O => \N__41327\,
            I => \N__41320\
        );

    \I__9418\ : InMux
    port map (
            O => \N__41326\,
            I => \N__41320\
        );

    \I__9417\ : InMux
    port map (
            O => \N__41325\,
            I => \N__41317\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__41320\,
            I => \N__41314\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__41317\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__9414\ : Odrv4
    port map (
            O => \N__41314\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__9413\ : InMux
    port map (
            O => \N__41309\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__9412\ : InMux
    port map (
            O => \N__41306\,
            I => \N__41303\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__41303\,
            I => \N__41299\
        );

    \I__9410\ : InMux
    port map (
            O => \N__41302\,
            I => \N__41296\
        );

    \I__9409\ : Span4Mux_h
    port map (
            O => \N__41299\,
            I => \N__41293\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__41296\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__9407\ : Odrv4
    port map (
            O => \N__41293\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__9406\ : InMux
    port map (
            O => \N__41288\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__9405\ : CascadeMux
    port map (
            O => \N__41285\,
            I => \N__41282\
        );

    \I__9404\ : InMux
    port map (
            O => \N__41282\,
            I => \N__41278\
        );

    \I__9403\ : InMux
    port map (
            O => \N__41281\,
            I => \N__41274\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__41278\,
            I => \N__41271\
        );

    \I__9401\ : InMux
    port map (
            O => \N__41277\,
            I => \N__41268\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__41274\,
            I => \N__41263\
        );

    \I__9399\ : Span4Mux_h
    port map (
            O => \N__41271\,
            I => \N__41263\
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__41268\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__9397\ : Odrv4
    port map (
            O => \N__41263\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__9396\ : InMux
    port map (
            O => \N__41258\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__9395\ : InMux
    port map (
            O => \N__41255\,
            I => \N__41248\
        );

    \I__9394\ : InMux
    port map (
            O => \N__41254\,
            I => \N__41248\
        );

    \I__9393\ : InMux
    port map (
            O => \N__41253\,
            I => \N__41245\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__41248\,
            I => \N__41242\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__41245\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__9390\ : Odrv4
    port map (
            O => \N__41242\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__9389\ : InMux
    port map (
            O => \N__41237\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__9388\ : CascadeMux
    port map (
            O => \N__41234\,
            I => \N__41230\
        );

    \I__9387\ : CascadeMux
    port map (
            O => \N__41233\,
            I => \N__41227\
        );

    \I__9386\ : InMux
    port map (
            O => \N__41230\,
            I => \N__41221\
        );

    \I__9385\ : InMux
    port map (
            O => \N__41227\,
            I => \N__41221\
        );

    \I__9384\ : InMux
    port map (
            O => \N__41226\,
            I => \N__41218\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__41221\,
            I => \N__41215\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__41218\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__9381\ : Odrv4
    port map (
            O => \N__41215\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__9380\ : InMux
    port map (
            O => \N__41210\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__9379\ : InMux
    port map (
            O => \N__41207\,
            I => \N__41203\
        );

    \I__9378\ : CascadeMux
    port map (
            O => \N__41206\,
            I => \N__41200\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__41203\,
            I => \N__41196\
        );

    \I__9376\ : InMux
    port map (
            O => \N__41200\,
            I => \N__41193\
        );

    \I__9375\ : InMux
    port map (
            O => \N__41199\,
            I => \N__41190\
        );

    \I__9374\ : Span4Mux_v
    port map (
            O => \N__41196\,
            I => \N__41185\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__41193\,
            I => \N__41185\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__41190\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__9371\ : Odrv4
    port map (
            O => \N__41185\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__9370\ : InMux
    port map (
            O => \N__41180\,
            I => \bfn_18_9_0_\
        );

    \I__9369\ : CascadeMux
    port map (
            O => \N__41177\,
            I => \N__41174\
        );

    \I__9368\ : InMux
    port map (
            O => \N__41174\,
            I => \N__41171\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__41171\,
            I => \N__41166\
        );

    \I__9366\ : InMux
    port map (
            O => \N__41170\,
            I => \N__41163\
        );

    \I__9365\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41160\
        );

    \I__9364\ : Span4Mux_v
    port map (
            O => \N__41166\,
            I => \N__41157\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__41163\,
            I => \N__41154\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__41160\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__9361\ : Odrv4
    port map (
            O => \N__41157\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__9360\ : Odrv4
    port map (
            O => \N__41154\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__9359\ : InMux
    port map (
            O => \N__41147\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__9358\ : CascadeMux
    port map (
            O => \N__41144\,
            I => \N__41140\
        );

    \I__9357\ : CascadeMux
    port map (
            O => \N__41143\,
            I => \N__41137\
        );

    \I__9356\ : InMux
    port map (
            O => \N__41140\,
            I => \N__41131\
        );

    \I__9355\ : InMux
    port map (
            O => \N__41137\,
            I => \N__41131\
        );

    \I__9354\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41128\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__41131\,
            I => \N__41125\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__41128\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__9351\ : Odrv4
    port map (
            O => \N__41125\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__9350\ : InMux
    port map (
            O => \N__41120\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__9349\ : InMux
    port map (
            O => \N__41117\,
            I => \N__41110\
        );

    \I__9348\ : InMux
    port map (
            O => \N__41116\,
            I => \N__41110\
        );

    \I__9347\ : InMux
    port map (
            O => \N__41115\,
            I => \N__41107\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__41110\,
            I => \N__41104\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__41107\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__9344\ : Odrv4
    port map (
            O => \N__41104\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__9343\ : InMux
    port map (
            O => \N__41099\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__9342\ : CascadeMux
    port map (
            O => \N__41096\,
            I => \N__41092\
        );

    \I__9341\ : InMux
    port map (
            O => \N__41095\,
            I => \N__41089\
        );

    \I__9340\ : InMux
    port map (
            O => \N__41092\,
            I => \N__41085\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__41089\,
            I => \N__41082\
        );

    \I__9338\ : InMux
    port map (
            O => \N__41088\,
            I => \N__41079\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__41085\,
            I => \N__41074\
        );

    \I__9336\ : Span4Mux_h
    port map (
            O => \N__41082\,
            I => \N__41074\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__41079\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__9334\ : Odrv4
    port map (
            O => \N__41074\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__9333\ : InMux
    port map (
            O => \N__41069\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__9332\ : CascadeMux
    port map (
            O => \N__41066\,
            I => \N__41062\
        );

    \I__9331\ : InMux
    port map (
            O => \N__41065\,
            I => \N__41059\
        );

    \I__9330\ : InMux
    port map (
            O => \N__41062\,
            I => \N__41055\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__41059\,
            I => \N__41052\
        );

    \I__9328\ : InMux
    port map (
            O => \N__41058\,
            I => \N__41049\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__41055\,
            I => \N__41044\
        );

    \I__9326\ : Span4Mux_h
    port map (
            O => \N__41052\,
            I => \N__41044\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__41049\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__9324\ : Odrv4
    port map (
            O => \N__41044\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__9323\ : InMux
    port map (
            O => \N__41039\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__9322\ : CascadeMux
    port map (
            O => \N__41036\,
            I => \N__41033\
        );

    \I__9321\ : InMux
    port map (
            O => \N__41033\,
            I => \N__41029\
        );

    \I__9320\ : InMux
    port map (
            O => \N__41032\,
            I => \N__41025\
        );

    \I__9319\ : LocalMux
    port map (
            O => \N__41029\,
            I => \N__41022\
        );

    \I__9318\ : InMux
    port map (
            O => \N__41028\,
            I => \N__41019\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__41025\,
            I => \N__41014\
        );

    \I__9316\ : Span4Mux_h
    port map (
            O => \N__41022\,
            I => \N__41014\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__41019\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__9314\ : Odrv4
    port map (
            O => \N__41014\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__9313\ : InMux
    port map (
            O => \N__41009\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__9312\ : InMux
    port map (
            O => \N__41006\,
            I => \N__40999\
        );

    \I__9311\ : InMux
    port map (
            O => \N__41005\,
            I => \N__40999\
        );

    \I__9310\ : InMux
    port map (
            O => \N__41004\,
            I => \N__40996\
        );

    \I__9309\ : LocalMux
    port map (
            O => \N__40999\,
            I => \N__40993\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__40996\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__9307\ : Odrv4
    port map (
            O => \N__40993\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__9306\ : InMux
    port map (
            O => \N__40988\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__9305\ : CascadeMux
    port map (
            O => \N__40985\,
            I => \N__40981\
        );

    \I__9304\ : CascadeMux
    port map (
            O => \N__40984\,
            I => \N__40978\
        );

    \I__9303\ : InMux
    port map (
            O => \N__40981\,
            I => \N__40972\
        );

    \I__9302\ : InMux
    port map (
            O => \N__40978\,
            I => \N__40972\
        );

    \I__9301\ : InMux
    port map (
            O => \N__40977\,
            I => \N__40969\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__40972\,
            I => \N__40966\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__40969\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__9298\ : Odrv4
    port map (
            O => \N__40966\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__9297\ : InMux
    port map (
            O => \N__40961\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__9296\ : InMux
    port map (
            O => \N__40958\,
            I => \N__40954\
        );

    \I__9295\ : CascadeMux
    port map (
            O => \N__40957\,
            I => \N__40951\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__40954\,
            I => \N__40947\
        );

    \I__9293\ : InMux
    port map (
            O => \N__40951\,
            I => \N__40944\
        );

    \I__9292\ : InMux
    port map (
            O => \N__40950\,
            I => \N__40941\
        );

    \I__9291\ : Span4Mux_v
    port map (
            O => \N__40947\,
            I => \N__40936\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__40944\,
            I => \N__40936\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__40941\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__9288\ : Odrv4
    port map (
            O => \N__40936\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__9287\ : InMux
    port map (
            O => \N__40931\,
            I => \bfn_18_8_0_\
        );

    \I__9286\ : CascadeMux
    port map (
            O => \N__40928\,
            I => \N__40925\
        );

    \I__9285\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40921\
        );

    \I__9284\ : InMux
    port map (
            O => \N__40924\,
            I => \N__40917\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__40921\,
            I => \N__40914\
        );

    \I__9282\ : InMux
    port map (
            O => \N__40920\,
            I => \N__40911\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__40917\,
            I => \N__40906\
        );

    \I__9280\ : Span4Mux_v
    port map (
            O => \N__40914\,
            I => \N__40906\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__40911\,
            I => \N__40903\
        );

    \I__9278\ : Odrv4
    port map (
            O => \N__40906\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__9277\ : Odrv4
    port map (
            O => \N__40903\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__9276\ : InMux
    port map (
            O => \N__40898\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__9275\ : CascadeMux
    port map (
            O => \N__40895\,
            I => \N__40891\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__40894\,
            I => \N__40888\
        );

    \I__9273\ : InMux
    port map (
            O => \N__40891\,
            I => \N__40882\
        );

    \I__9272\ : InMux
    port map (
            O => \N__40888\,
            I => \N__40882\
        );

    \I__9271\ : InMux
    port map (
            O => \N__40887\,
            I => \N__40879\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__40882\,
            I => \N__40876\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__40879\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__9268\ : Odrv4
    port map (
            O => \N__40876\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__9267\ : InMux
    port map (
            O => \N__40871\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__9266\ : InMux
    port map (
            O => \N__40868\,
            I => \N__40861\
        );

    \I__9265\ : InMux
    port map (
            O => \N__40867\,
            I => \N__40861\
        );

    \I__9264\ : InMux
    port map (
            O => \N__40866\,
            I => \N__40858\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__40861\,
            I => \N__40855\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__40858\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__9261\ : Odrv4
    port map (
            O => \N__40855\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__9260\ : InMux
    port map (
            O => \N__40850\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__9259\ : CascadeMux
    port map (
            O => \N__40847\,
            I => \N__40843\
        );

    \I__9258\ : InMux
    port map (
            O => \N__40846\,
            I => \N__40840\
        );

    \I__9257\ : InMux
    port map (
            O => \N__40843\,
            I => \N__40836\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__40840\,
            I => \N__40833\
        );

    \I__9255\ : InMux
    port map (
            O => \N__40839\,
            I => \N__40830\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__40836\,
            I => \N__40825\
        );

    \I__9253\ : Span4Mux_h
    port map (
            O => \N__40833\,
            I => \N__40825\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__40830\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__9251\ : Odrv4
    port map (
            O => \N__40825\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__9250\ : InMux
    port map (
            O => \N__40820\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__9249\ : CascadeMux
    port map (
            O => \N__40817\,
            I => \phase_controller_inst2.stoper_tr.N_45_cascade_\
        );

    \I__9248\ : InMux
    port map (
            O => \N__40814\,
            I => \N__40810\
        );

    \I__9247\ : InMux
    port map (
            O => \N__40813\,
            I => \N__40807\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__40810\,
            I => \N__40804\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__40807\,
            I => \N__40801\
        );

    \I__9244\ : Span4Mux_h
    port map (
            O => \N__40804\,
            I => \N__40797\
        );

    \I__9243\ : Span4Mux_v
    port map (
            O => \N__40801\,
            I => \N__40794\
        );

    \I__9242\ : InMux
    port map (
            O => \N__40800\,
            I => \N__40791\
        );

    \I__9241\ : Span4Mux_h
    port map (
            O => \N__40797\,
            I => \N__40788\
        );

    \I__9240\ : Span4Mux_h
    port map (
            O => \N__40794\,
            I => \N__40785\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__40791\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__9238\ : Odrv4
    port map (
            O => \N__40788\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__9237\ : Odrv4
    port map (
            O => \N__40785\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__9236\ : InMux
    port map (
            O => \N__40778\,
            I => \N__40774\
        );

    \I__9235\ : InMux
    port map (
            O => \N__40777\,
            I => \N__40771\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__40774\,
            I => \N__40766\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__40771\,
            I => \N__40766\
        );

    \I__9232\ : Span4Mux_v
    port map (
            O => \N__40766\,
            I => \N__40762\
        );

    \I__9231\ : InMux
    port map (
            O => \N__40765\,
            I => \N__40759\
        );

    \I__9230\ : Odrv4
    port map (
            O => \N__40762\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__40759\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__9228\ : InMux
    port map (
            O => \N__40754\,
            I => \bfn_18_7_0_\
        );

    \I__9227\ : CascadeMux
    port map (
            O => \N__40751\,
            I => \N__40747\
        );

    \I__9226\ : InMux
    port map (
            O => \N__40750\,
            I => \N__40744\
        );

    \I__9225\ : InMux
    port map (
            O => \N__40747\,
            I => \N__40741\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__40744\,
            I => \N__40735\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__40741\,
            I => \N__40735\
        );

    \I__9222\ : InMux
    port map (
            O => \N__40740\,
            I => \N__40732\
        );

    \I__9221\ : Span4Mux_v
    port map (
            O => \N__40735\,
            I => \N__40729\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__40732\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__9219\ : Odrv4
    port map (
            O => \N__40729\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__9218\ : InMux
    port map (
            O => \N__40724\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__9217\ : CascadeMux
    port map (
            O => \N__40721\,
            I => \N__40717\
        );

    \I__9216\ : CascadeMux
    port map (
            O => \N__40720\,
            I => \N__40714\
        );

    \I__9215\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40708\
        );

    \I__9214\ : InMux
    port map (
            O => \N__40714\,
            I => \N__40708\
        );

    \I__9213\ : InMux
    port map (
            O => \N__40713\,
            I => \N__40705\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__40708\,
            I => \N__40702\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__40705\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__9210\ : Odrv4
    port map (
            O => \N__40702\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__9209\ : InMux
    port map (
            O => \N__40697\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__9208\ : InMux
    port map (
            O => \N__40694\,
            I => \N__40687\
        );

    \I__9207\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40687\
        );

    \I__9206\ : InMux
    port map (
            O => \N__40692\,
            I => \N__40684\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__40687\,
            I => \N__40681\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__40684\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__9203\ : Odrv4
    port map (
            O => \N__40681\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__9202\ : InMux
    port map (
            O => \N__40676\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__9201\ : CascadeMux
    port map (
            O => \N__40673\,
            I => \N__40670\
        );

    \I__9200\ : InMux
    port map (
            O => \N__40670\,
            I => \N__40667\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__40667\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__9198\ : InMux
    port map (
            O => \N__40664\,
            I => \N__40661\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__40661\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__9196\ : CascadeMux
    port map (
            O => \N__40658\,
            I => \N__40655\
        );

    \I__9195\ : InMux
    port map (
            O => \N__40655\,
            I => \N__40652\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__40652\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__9193\ : InMux
    port map (
            O => \N__40649\,
            I => \N__40646\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__40646\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__9191\ : CascadeMux
    port map (
            O => \N__40643\,
            I => \N__40640\
        );

    \I__9190\ : InMux
    port map (
            O => \N__40640\,
            I => \N__40637\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__40637\,
            I => \N__40634\
        );

    \I__9188\ : Span4Mux_h
    port map (
            O => \N__40634\,
            I => \N__40631\
        );

    \I__9187\ : Odrv4
    port map (
            O => \N__40631\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__9186\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40625\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__40625\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__9184\ : CascadeMux
    port map (
            O => \N__40622\,
            I => \N__40603\
        );

    \I__9183\ : CascadeMux
    port map (
            O => \N__40621\,
            I => \N__40599\
        );

    \I__9182\ : CascadeMux
    port map (
            O => \N__40620\,
            I => \N__40595\
        );

    \I__9181\ : CascadeMux
    port map (
            O => \N__40619\,
            I => \N__40591\
        );

    \I__9180\ : CascadeMux
    port map (
            O => \N__40618\,
            I => \N__40587\
        );

    \I__9179\ : CascadeMux
    port map (
            O => \N__40617\,
            I => \N__40583\
        );

    \I__9178\ : CascadeMux
    port map (
            O => \N__40616\,
            I => \N__40579\
        );

    \I__9177\ : InMux
    port map (
            O => \N__40615\,
            I => \N__40564\
        );

    \I__9176\ : InMux
    port map (
            O => \N__40614\,
            I => \N__40564\
        );

    \I__9175\ : InMux
    port map (
            O => \N__40613\,
            I => \N__40564\
        );

    \I__9174\ : InMux
    port map (
            O => \N__40612\,
            I => \N__40561\
        );

    \I__9173\ : InMux
    port map (
            O => \N__40611\,
            I => \N__40552\
        );

    \I__9172\ : InMux
    port map (
            O => \N__40610\,
            I => \N__40552\
        );

    \I__9171\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40552\
        );

    \I__9170\ : InMux
    port map (
            O => \N__40608\,
            I => \N__40552\
        );

    \I__9169\ : CascadeMux
    port map (
            O => \N__40607\,
            I => \N__40548\
        );

    \I__9168\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40532\
        );

    \I__9167\ : InMux
    port map (
            O => \N__40603\,
            I => \N__40532\
        );

    \I__9166\ : InMux
    port map (
            O => \N__40602\,
            I => \N__40532\
        );

    \I__9165\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40532\
        );

    \I__9164\ : InMux
    port map (
            O => \N__40598\,
            I => \N__40532\
        );

    \I__9163\ : InMux
    port map (
            O => \N__40595\,
            I => \N__40532\
        );

    \I__9162\ : InMux
    port map (
            O => \N__40594\,
            I => \N__40532\
        );

    \I__9161\ : InMux
    port map (
            O => \N__40591\,
            I => \N__40515\
        );

    \I__9160\ : InMux
    port map (
            O => \N__40590\,
            I => \N__40515\
        );

    \I__9159\ : InMux
    port map (
            O => \N__40587\,
            I => \N__40515\
        );

    \I__9158\ : InMux
    port map (
            O => \N__40586\,
            I => \N__40515\
        );

    \I__9157\ : InMux
    port map (
            O => \N__40583\,
            I => \N__40515\
        );

    \I__9156\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40515\
        );

    \I__9155\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40515\
        );

    \I__9154\ : InMux
    port map (
            O => \N__40578\,
            I => \N__40515\
        );

    \I__9153\ : CascadeMux
    port map (
            O => \N__40577\,
            I => \N__40511\
        );

    \I__9152\ : CascadeMux
    port map (
            O => \N__40576\,
            I => \N__40507\
        );

    \I__9151\ : CascadeMux
    port map (
            O => \N__40575\,
            I => \N__40503\
        );

    \I__9150\ : CascadeMux
    port map (
            O => \N__40574\,
            I => \N__40499\
        );

    \I__9149\ : CascadeMux
    port map (
            O => \N__40573\,
            I => \N__40495\
        );

    \I__9148\ : CascadeMux
    port map (
            O => \N__40572\,
            I => \N__40491\
        );

    \I__9147\ : CascadeMux
    port map (
            O => \N__40571\,
            I => \N__40487\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__40564\,
            I => \N__40482\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__40561\,
            I => \N__40477\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__40552\,
            I => \N__40477\
        );

    \I__9143\ : InMux
    port map (
            O => \N__40551\,
            I => \N__40470\
        );

    \I__9142\ : InMux
    port map (
            O => \N__40548\,
            I => \N__40470\
        );

    \I__9141\ : InMux
    port map (
            O => \N__40547\,
            I => \N__40470\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__40532\,
            I => \N__40458\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__40515\,
            I => \N__40455\
        );

    \I__9138\ : InMux
    port map (
            O => \N__40514\,
            I => \N__40438\
        );

    \I__9137\ : InMux
    port map (
            O => \N__40511\,
            I => \N__40438\
        );

    \I__9136\ : InMux
    port map (
            O => \N__40510\,
            I => \N__40438\
        );

    \I__9135\ : InMux
    port map (
            O => \N__40507\,
            I => \N__40438\
        );

    \I__9134\ : InMux
    port map (
            O => \N__40506\,
            I => \N__40438\
        );

    \I__9133\ : InMux
    port map (
            O => \N__40503\,
            I => \N__40438\
        );

    \I__9132\ : InMux
    port map (
            O => \N__40502\,
            I => \N__40438\
        );

    \I__9131\ : InMux
    port map (
            O => \N__40499\,
            I => \N__40438\
        );

    \I__9130\ : InMux
    port map (
            O => \N__40498\,
            I => \N__40423\
        );

    \I__9129\ : InMux
    port map (
            O => \N__40495\,
            I => \N__40423\
        );

    \I__9128\ : InMux
    port map (
            O => \N__40494\,
            I => \N__40423\
        );

    \I__9127\ : InMux
    port map (
            O => \N__40491\,
            I => \N__40423\
        );

    \I__9126\ : InMux
    port map (
            O => \N__40490\,
            I => \N__40423\
        );

    \I__9125\ : InMux
    port map (
            O => \N__40487\,
            I => \N__40423\
        );

    \I__9124\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40423\
        );

    \I__9123\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40420\
        );

    \I__9122\ : Span4Mux_v
    port map (
            O => \N__40482\,
            I => \N__40413\
        );

    \I__9121\ : Span4Mux_v
    port map (
            O => \N__40477\,
            I => \N__40413\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__40470\,
            I => \N__40413\
        );

    \I__9119\ : InMux
    port map (
            O => \N__40469\,
            I => \N__40410\
        );

    \I__9118\ : InMux
    port map (
            O => \N__40468\,
            I => \N__40403\
        );

    \I__9117\ : InMux
    port map (
            O => \N__40467\,
            I => \N__40403\
        );

    \I__9116\ : InMux
    port map (
            O => \N__40466\,
            I => \N__40403\
        );

    \I__9115\ : InMux
    port map (
            O => \N__40465\,
            I => \N__40394\
        );

    \I__9114\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40394\
        );

    \I__9113\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40394\
        );

    \I__9112\ : InMux
    port map (
            O => \N__40462\,
            I => \N__40394\
        );

    \I__9111\ : InMux
    port map (
            O => \N__40461\,
            I => \N__40391\
        );

    \I__9110\ : Span4Mux_v
    port map (
            O => \N__40458\,
            I => \N__40382\
        );

    \I__9109\ : Span4Mux_h
    port map (
            O => \N__40455\,
            I => \N__40382\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__40438\,
            I => \N__40382\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__40423\,
            I => \N__40382\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__40420\,
            I => \N__40379\
        );

    \I__9105\ : Span4Mux_v
    port map (
            O => \N__40413\,
            I => \N__40373\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__40410\,
            I => \N__40366\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__40403\,
            I => \N__40366\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__40394\,
            I => \N__40366\
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__40391\,
            I => \N__40363\
        );

    \I__9100\ : Span4Mux_v
    port map (
            O => \N__40382\,
            I => \N__40360\
        );

    \I__9099\ : Span4Mux_v
    port map (
            O => \N__40379\,
            I => \N__40357\
        );

    \I__9098\ : InMux
    port map (
            O => \N__40378\,
            I => \N__40354\
        );

    \I__9097\ : InMux
    port map (
            O => \N__40377\,
            I => \N__40351\
        );

    \I__9096\ : InMux
    port map (
            O => \N__40376\,
            I => \N__40348\
        );

    \I__9095\ : Span4Mux_v
    port map (
            O => \N__40373\,
            I => \N__40345\
        );

    \I__9094\ : Span4Mux_v
    port map (
            O => \N__40366\,
            I => \N__40342\
        );

    \I__9093\ : Sp12to4
    port map (
            O => \N__40363\,
            I => \N__40339\
        );

    \I__9092\ : Span4Mux_v
    port map (
            O => \N__40360\,
            I => \N__40336\
        );

    \I__9091\ : Sp12to4
    port map (
            O => \N__40357\,
            I => \N__40333\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__40354\,
            I => \N__40326\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__40351\,
            I => \N__40326\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__40348\,
            I => \N__40326\
        );

    \I__9087\ : Span4Mux_v
    port map (
            O => \N__40345\,
            I => \N__40323\
        );

    \I__9086\ : Span4Mux_h
    port map (
            O => \N__40342\,
            I => \N__40320\
        );

    \I__9085\ : Span12Mux_v
    port map (
            O => \N__40339\,
            I => \N__40313\
        );

    \I__9084\ : Sp12to4
    port map (
            O => \N__40336\,
            I => \N__40313\
        );

    \I__9083\ : Span12Mux_s9_h
    port map (
            O => \N__40333\,
            I => \N__40313\
        );

    \I__9082\ : IoSpan4Mux
    port map (
            O => \N__40326\,
            I => \N__40310\
        );

    \I__9081\ : Span4Mux_v
    port map (
            O => \N__40323\,
            I => \N__40307\
        );

    \I__9080\ : Sp12to4
    port map (
            O => \N__40320\,
            I => \N__40302\
        );

    \I__9079\ : Span12Mux_h
    port map (
            O => \N__40313\,
            I => \N__40302\
        );

    \I__9078\ : Span4Mux_s3_v
    port map (
            O => \N__40310\,
            I => \N__40299\
        );

    \I__9077\ : Odrv4
    port map (
            O => \N__40307\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9076\ : Odrv12
    port map (
            O => \N__40302\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9075\ : Odrv4
    port map (
            O => \N__40299\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9074\ : CascadeMux
    port map (
            O => \N__40292\,
            I => \N__40289\
        );

    \I__9073\ : InMux
    port map (
            O => \N__40289\,
            I => \N__40286\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__40286\,
            I => \N__40283\
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__40283\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__9070\ : CascadeMux
    port map (
            O => \N__40280\,
            I => \N__40266\
        );

    \I__9069\ : CascadeMux
    port map (
            O => \N__40279\,
            I => \N__40262\
        );

    \I__9068\ : CascadeMux
    port map (
            O => \N__40278\,
            I => \N__40259\
        );

    \I__9067\ : CascadeMux
    port map (
            O => \N__40277\,
            I => \N__40256\
        );

    \I__9066\ : CascadeMux
    port map (
            O => \N__40276\,
            I => \N__40252\
        );

    \I__9065\ : CascadeMux
    port map (
            O => \N__40275\,
            I => \N__40249\
        );

    \I__9064\ : CascadeMux
    port map (
            O => \N__40274\,
            I => \N__40245\
        );

    \I__9063\ : CascadeMux
    port map (
            O => \N__40273\,
            I => \N__40242\
        );

    \I__9062\ : CascadeMux
    port map (
            O => \N__40272\,
            I => \N__40239\
        );

    \I__9061\ : CascadeMux
    port map (
            O => \N__40271\,
            I => \N__40236\
        );

    \I__9060\ : CascadeMux
    port map (
            O => \N__40270\,
            I => \N__40233\
        );

    \I__9059\ : CascadeMux
    port map (
            O => \N__40269\,
            I => \N__40230\
        );

    \I__9058\ : InMux
    port map (
            O => \N__40266\,
            I => \N__40207\
        );

    \I__9057\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40207\
        );

    \I__9056\ : InMux
    port map (
            O => \N__40262\,
            I => \N__40207\
        );

    \I__9055\ : InMux
    port map (
            O => \N__40259\,
            I => \N__40207\
        );

    \I__9054\ : InMux
    port map (
            O => \N__40256\,
            I => \N__40207\
        );

    \I__9053\ : InMux
    port map (
            O => \N__40255\,
            I => \N__40194\
        );

    \I__9052\ : InMux
    port map (
            O => \N__40252\,
            I => \N__40194\
        );

    \I__9051\ : InMux
    port map (
            O => \N__40249\,
            I => \N__40194\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40248\,
            I => \N__40194\
        );

    \I__9049\ : InMux
    port map (
            O => \N__40245\,
            I => \N__40194\
        );

    \I__9048\ : InMux
    port map (
            O => \N__40242\,
            I => \N__40194\
        );

    \I__9047\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40185\
        );

    \I__9046\ : InMux
    port map (
            O => \N__40236\,
            I => \N__40185\
        );

    \I__9045\ : InMux
    port map (
            O => \N__40233\,
            I => \N__40185\
        );

    \I__9044\ : InMux
    port map (
            O => \N__40230\,
            I => \N__40185\
        );

    \I__9043\ : CascadeMux
    port map (
            O => \N__40229\,
            I => \N__40178\
        );

    \I__9042\ : CascadeMux
    port map (
            O => \N__40228\,
            I => \N__40175\
        );

    \I__9041\ : CascadeMux
    port map (
            O => \N__40227\,
            I => \N__40172\
        );

    \I__9040\ : CascadeMux
    port map (
            O => \N__40226\,
            I => \N__40169\
        );

    \I__9039\ : CascadeMux
    port map (
            O => \N__40225\,
            I => \N__40165\
        );

    \I__9038\ : CascadeMux
    port map (
            O => \N__40224\,
            I => \N__40161\
        );

    \I__9037\ : CascadeMux
    port map (
            O => \N__40223\,
            I => \N__40157\
        );

    \I__9036\ : CascadeMux
    port map (
            O => \N__40222\,
            I => \N__40153\
        );

    \I__9035\ : CascadeMux
    port map (
            O => \N__40221\,
            I => \N__40150\
        );

    \I__9034\ : CascadeMux
    port map (
            O => \N__40220\,
            I => \N__40147\
        );

    \I__9033\ : CascadeMux
    port map (
            O => \N__40219\,
            I => \N__40144\
        );

    \I__9032\ : InMux
    port map (
            O => \N__40218\,
            I => \N__40140\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__40207\,
            I => \N__40133\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__40194\,
            I => \N__40133\
        );

    \I__9029\ : LocalMux
    port map (
            O => \N__40185\,
            I => \N__40133\
        );

    \I__9028\ : InMux
    port map (
            O => \N__40184\,
            I => \N__40126\
        );

    \I__9027\ : InMux
    port map (
            O => \N__40183\,
            I => \N__40126\
        );

    \I__9026\ : InMux
    port map (
            O => \N__40182\,
            I => \N__40126\
        );

    \I__9025\ : InMux
    port map (
            O => \N__40181\,
            I => \N__40111\
        );

    \I__9024\ : InMux
    port map (
            O => \N__40178\,
            I => \N__40102\
        );

    \I__9023\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40102\
        );

    \I__9022\ : InMux
    port map (
            O => \N__40172\,
            I => \N__40097\
        );

    \I__9021\ : InMux
    port map (
            O => \N__40169\,
            I => \N__40097\
        );

    \I__9020\ : InMux
    port map (
            O => \N__40168\,
            I => \N__40080\
        );

    \I__9019\ : InMux
    port map (
            O => \N__40165\,
            I => \N__40080\
        );

    \I__9018\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40080\
        );

    \I__9017\ : InMux
    port map (
            O => \N__40161\,
            I => \N__40080\
        );

    \I__9016\ : InMux
    port map (
            O => \N__40160\,
            I => \N__40080\
        );

    \I__9015\ : InMux
    port map (
            O => \N__40157\,
            I => \N__40080\
        );

    \I__9014\ : InMux
    port map (
            O => \N__40156\,
            I => \N__40080\
        );

    \I__9013\ : InMux
    port map (
            O => \N__40153\,
            I => \N__40080\
        );

    \I__9012\ : InMux
    port map (
            O => \N__40150\,
            I => \N__40071\
        );

    \I__9011\ : InMux
    port map (
            O => \N__40147\,
            I => \N__40071\
        );

    \I__9010\ : InMux
    port map (
            O => \N__40144\,
            I => \N__40071\
        );

    \I__9009\ : InMux
    port map (
            O => \N__40143\,
            I => \N__40071\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__40140\,
            I => \N__40064\
        );

    \I__9007\ : Span4Mux_v
    port map (
            O => \N__40133\,
            I => \N__40064\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__40126\,
            I => \N__40064\
        );

    \I__9005\ : InMux
    port map (
            O => \N__40125\,
            I => \N__40058\
        );

    \I__9004\ : InMux
    port map (
            O => \N__40124\,
            I => \N__40052\
        );

    \I__9003\ : InMux
    port map (
            O => \N__40123\,
            I => \N__40052\
        );

    \I__9002\ : InMux
    port map (
            O => \N__40122\,
            I => \N__40037\
        );

    \I__9001\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40037\
        );

    \I__9000\ : InMux
    port map (
            O => \N__40120\,
            I => \N__40037\
        );

    \I__8999\ : InMux
    port map (
            O => \N__40119\,
            I => \N__40037\
        );

    \I__8998\ : InMux
    port map (
            O => \N__40118\,
            I => \N__40037\
        );

    \I__8997\ : InMux
    port map (
            O => \N__40117\,
            I => \N__40037\
        );

    \I__8996\ : InMux
    port map (
            O => \N__40116\,
            I => \N__40037\
        );

    \I__8995\ : InMux
    port map (
            O => \N__40115\,
            I => \N__40032\
        );

    \I__8994\ : InMux
    port map (
            O => \N__40114\,
            I => \N__40032\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__40111\,
            I => \N__40029\
        );

    \I__8992\ : InMux
    port map (
            O => \N__40110\,
            I => \N__40020\
        );

    \I__8991\ : InMux
    port map (
            O => \N__40109\,
            I => \N__40020\
        );

    \I__8990\ : InMux
    port map (
            O => \N__40108\,
            I => \N__40020\
        );

    \I__8989\ : InMux
    port map (
            O => \N__40107\,
            I => \N__40020\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__40102\,
            I => \N__40009\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__40097\,
            I => \N__40009\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__40080\,
            I => \N__40009\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__40071\,
            I => \N__40009\
        );

    \I__8984\ : Span4Mux_h
    port map (
            O => \N__40064\,
            I => \N__40009\
        );

    \I__8983\ : InMux
    port map (
            O => \N__40063\,
            I => \N__40004\
        );

    \I__8982\ : InMux
    port map (
            O => \N__40062\,
            I => \N__40004\
        );

    \I__8981\ : InMux
    port map (
            O => \N__40061\,
            I => \N__40000\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__40058\,
            I => \N__39992\
        );

    \I__8979\ : InMux
    port map (
            O => \N__40057\,
            I => \N__39988\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__40052\,
            I => \N__39981\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__40037\,
            I => \N__39981\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__40032\,
            I => \N__39981\
        );

    \I__8975\ : Span4Mux_v
    port map (
            O => \N__40029\,
            I => \N__39964\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__40020\,
            I => \N__39964\
        );

    \I__8973\ : Span4Mux_v
    port map (
            O => \N__40009\,
            I => \N__39964\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__40004\,
            I => \N__39964\
        );

    \I__8971\ : InMux
    port map (
            O => \N__40003\,
            I => \N__39954\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__40000\,
            I => \N__39951\
        );

    \I__8969\ : InMux
    port map (
            O => \N__39999\,
            I => \N__39940\
        );

    \I__8968\ : InMux
    port map (
            O => \N__39998\,
            I => \N__39940\
        );

    \I__8967\ : InMux
    port map (
            O => \N__39997\,
            I => \N__39940\
        );

    \I__8966\ : InMux
    port map (
            O => \N__39996\,
            I => \N__39940\
        );

    \I__8965\ : InMux
    port map (
            O => \N__39995\,
            I => \N__39940\
        );

    \I__8964\ : Span12Mux_s11_v
    port map (
            O => \N__39992\,
            I => \N__39937\
        );

    \I__8963\ : InMux
    port map (
            O => \N__39991\,
            I => \N__39934\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__39988\,
            I => \N__39929\
        );

    \I__8961\ : Span4Mux_v
    port map (
            O => \N__39981\,
            I => \N__39929\
        );

    \I__8960\ : InMux
    port map (
            O => \N__39980\,
            I => \N__39926\
        );

    \I__8959\ : InMux
    port map (
            O => \N__39979\,
            I => \N__39911\
        );

    \I__8958\ : InMux
    port map (
            O => \N__39978\,
            I => \N__39911\
        );

    \I__8957\ : InMux
    port map (
            O => \N__39977\,
            I => \N__39911\
        );

    \I__8956\ : InMux
    port map (
            O => \N__39976\,
            I => \N__39911\
        );

    \I__8955\ : InMux
    port map (
            O => \N__39975\,
            I => \N__39911\
        );

    \I__8954\ : InMux
    port map (
            O => \N__39974\,
            I => \N__39911\
        );

    \I__8953\ : InMux
    port map (
            O => \N__39973\,
            I => \N__39911\
        );

    \I__8952\ : Span4Mux_h
    port map (
            O => \N__39964\,
            I => \N__39908\
        );

    \I__8951\ : InMux
    port map (
            O => \N__39963\,
            I => \N__39893\
        );

    \I__8950\ : InMux
    port map (
            O => \N__39962\,
            I => \N__39893\
        );

    \I__8949\ : InMux
    port map (
            O => \N__39961\,
            I => \N__39893\
        );

    \I__8948\ : InMux
    port map (
            O => \N__39960\,
            I => \N__39893\
        );

    \I__8947\ : InMux
    port map (
            O => \N__39959\,
            I => \N__39893\
        );

    \I__8946\ : InMux
    port map (
            O => \N__39958\,
            I => \N__39893\
        );

    \I__8945\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39893\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__39954\,
            I => \N__39886\
        );

    \I__8943\ : Span12Mux_h
    port map (
            O => \N__39951\,
            I => \N__39886\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__39940\,
            I => \N__39886\
        );

    \I__8941\ : Odrv12
    port map (
            O => \N__39937\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__39934\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8939\ : Odrv4
    port map (
            O => \N__39929\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__39926\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__39911\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8936\ : Odrv4
    port map (
            O => \N__39908\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__39893\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8934\ : Odrv12
    port map (
            O => \N__39886\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8933\ : InMux
    port map (
            O => \N__39869\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__8932\ : CascadeMux
    port map (
            O => \N__39866\,
            I => \N__39861\
        );

    \I__8931\ : CascadeMux
    port map (
            O => \N__39865\,
            I => \N__39858\
        );

    \I__8930\ : InMux
    port map (
            O => \N__39864\,
            I => \N__39854\
        );

    \I__8929\ : InMux
    port map (
            O => \N__39861\,
            I => \N__39851\
        );

    \I__8928\ : InMux
    port map (
            O => \N__39858\,
            I => \N__39848\
        );

    \I__8927\ : InMux
    port map (
            O => \N__39857\,
            I => \N__39845\
        );

    \I__8926\ : LocalMux
    port map (
            O => \N__39854\,
            I => \N__39842\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__39851\,
            I => \N__39839\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__39848\,
            I => \N__39836\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__39845\,
            I => \N__39833\
        );

    \I__8922\ : Span4Mux_h
    port map (
            O => \N__39842\,
            I => \N__39828\
        );

    \I__8921\ : Span4Mux_h
    port map (
            O => \N__39839\,
            I => \N__39828\
        );

    \I__8920\ : Span4Mux_h
    port map (
            O => \N__39836\,
            I => \N__39825\
        );

    \I__8919\ : Span12Mux_v
    port map (
            O => \N__39833\,
            I => \N__39822\
        );

    \I__8918\ : Span4Mux_h
    port map (
            O => \N__39828\,
            I => \N__39819\
        );

    \I__8917\ : Span4Mux_h
    port map (
            O => \N__39825\,
            I => \N__39816\
        );

    \I__8916\ : Odrv12
    port map (
            O => \N__39822\,
            I => \current_shift_inst.N_1310_i\
        );

    \I__8915\ : Odrv4
    port map (
            O => \N__39819\,
            I => \current_shift_inst.N_1310_i\
        );

    \I__8914\ : Odrv4
    port map (
            O => \N__39816\,
            I => \current_shift_inst.N_1310_i\
        );

    \I__8913\ : InMux
    port map (
            O => \N__39809\,
            I => \N__39806\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__39806\,
            I => \N__39803\
        );

    \I__8911\ : Odrv4
    port map (
            O => \N__39803\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__8910\ : CascadeMux
    port map (
            O => \N__39800\,
            I => \N__39797\
        );

    \I__8909\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39794\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__39794\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__8907\ : InMux
    port map (
            O => \N__39791\,
            I => \N__39788\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__39788\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__8905\ : CascadeMux
    port map (
            O => \N__39785\,
            I => \N__39782\
        );

    \I__8904\ : InMux
    port map (
            O => \N__39782\,
            I => \N__39779\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__39779\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__8902\ : InMux
    port map (
            O => \N__39776\,
            I => \N__39773\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__39773\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__8900\ : CascadeMux
    port map (
            O => \N__39770\,
            I => \N__39767\
        );

    \I__8899\ : InMux
    port map (
            O => \N__39767\,
            I => \N__39764\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__39764\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__8897\ : InMux
    port map (
            O => \N__39761\,
            I => \N__39758\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__39758\,
            I => \N__39755\
        );

    \I__8895\ : Odrv4
    port map (
            O => \N__39755\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__8894\ : CascadeMux
    port map (
            O => \N__39752\,
            I => \N__39749\
        );

    \I__8893\ : InMux
    port map (
            O => \N__39749\,
            I => \N__39746\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__39746\,
            I => \N__39743\
        );

    \I__8891\ : Odrv4
    port map (
            O => \N__39743\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__8890\ : CascadeMux
    port map (
            O => \N__39740\,
            I => \N__39737\
        );

    \I__8889\ : InMux
    port map (
            O => \N__39737\,
            I => \N__39734\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__39734\,
            I => \N__39731\
        );

    \I__8887\ : Odrv4
    port map (
            O => \N__39731\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__8886\ : CascadeMux
    port map (
            O => \N__39728\,
            I => \N__39725\
        );

    \I__8885\ : InMux
    port map (
            O => \N__39725\,
            I => \N__39722\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__39722\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__8883\ : InMux
    port map (
            O => \N__39719\,
            I => \N__39716\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__39716\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__8881\ : CascadeMux
    port map (
            O => \N__39713\,
            I => \N__39710\
        );

    \I__8880\ : InMux
    port map (
            O => \N__39710\,
            I => \N__39707\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__39707\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__8878\ : InMux
    port map (
            O => \N__39704\,
            I => \N__39701\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__39701\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__8876\ : CascadeMux
    port map (
            O => \N__39698\,
            I => \N__39695\
        );

    \I__8875\ : InMux
    port map (
            O => \N__39695\,
            I => \N__39692\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__39692\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__8873\ : InMux
    port map (
            O => \N__39689\,
            I => \N__39686\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__39686\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__8871\ : CascadeMux
    port map (
            O => \N__39683\,
            I => \N__39680\
        );

    \I__8870\ : InMux
    port map (
            O => \N__39680\,
            I => \N__39677\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__39677\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__8868\ : InMux
    port map (
            O => \N__39674\,
            I => \N__39671\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__39671\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__8866\ : InMux
    port map (
            O => \N__39668\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__8865\ : SRMux
    port map (
            O => \N__39665\,
            I => \N__39661\
        );

    \I__8864\ : SRMux
    port map (
            O => \N__39664\,
            I => \N__39658\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__39661\,
            I => \N__39652\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__39658\,
            I => \N__39652\
        );

    \I__8861\ : SRMux
    port map (
            O => \N__39657\,
            I => \N__39648\
        );

    \I__8860\ : Span4Mux_v
    port map (
            O => \N__39652\,
            I => \N__39645\
        );

    \I__8859\ : SRMux
    port map (
            O => \N__39651\,
            I => \N__39642\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__39648\,
            I => \N__39639\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__39645\,
            I => \N__39634\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__39642\,
            I => \N__39634\
        );

    \I__8855\ : Span4Mux_h
    port map (
            O => \N__39639\,
            I => \N__39631\
        );

    \I__8854\ : Span4Mux_h
    port map (
            O => \N__39634\,
            I => \N__39628\
        );

    \I__8853\ : Odrv4
    port map (
            O => \N__39631\,
            I => \phase_controller_inst1.stoper_tr.un1_stoper_state12_1_0_i\
        );

    \I__8852\ : Odrv4
    port map (
            O => \N__39628\,
            I => \phase_controller_inst1.stoper_tr.un1_stoper_state12_1_0_i\
        );

    \I__8851\ : InMux
    port map (
            O => \N__39623\,
            I => \N__39620\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__39620\,
            I => \N__39617\
        );

    \I__8849\ : Span4Mux_h
    port map (
            O => \N__39617\,
            I => \N__39614\
        );

    \I__8848\ : Odrv4
    port map (
            O => \N__39614\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__8847\ : CascadeMux
    port map (
            O => \N__39611\,
            I => \N__39608\
        );

    \I__8846\ : InMux
    port map (
            O => \N__39608\,
            I => \N__39605\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__39605\,
            I => \N__39602\
        );

    \I__8844\ : Span4Mux_h
    port map (
            O => \N__39602\,
            I => \N__39599\
        );

    \I__8843\ : Odrv4
    port map (
            O => \N__39599\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__8842\ : CascadeMux
    port map (
            O => \N__39596\,
            I => \N__39593\
        );

    \I__8841\ : InMux
    port map (
            O => \N__39593\,
            I => \N__39590\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__39590\,
            I => \N__39587\
        );

    \I__8839\ : Span4Mux_v
    port map (
            O => \N__39587\,
            I => \N__39584\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__39584\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__8837\ : InMux
    port map (
            O => \N__39581\,
            I => \N__39578\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__39578\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__8835\ : CascadeMux
    port map (
            O => \N__39575\,
            I => \N__39572\
        );

    \I__8834\ : InMux
    port map (
            O => \N__39572\,
            I => \N__39569\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__39569\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__8832\ : InMux
    port map (
            O => \N__39566\,
            I => \N__39563\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__39563\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__8830\ : CascadeMux
    port map (
            O => \N__39560\,
            I => \N__39557\
        );

    \I__8829\ : InMux
    port map (
            O => \N__39557\,
            I => \N__39554\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__39554\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__8827\ : InMux
    port map (
            O => \N__39551\,
            I => \N__39548\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__39548\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__8825\ : InMux
    port map (
            O => \N__39545\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__8824\ : InMux
    port map (
            O => \N__39542\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__8823\ : InMux
    port map (
            O => \N__39539\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__8822\ : InMux
    port map (
            O => \N__39536\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__8821\ : InMux
    port map (
            O => \N__39533\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__8820\ : InMux
    port map (
            O => \N__39530\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__8819\ : InMux
    port map (
            O => \N__39527\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__8818\ : InMux
    port map (
            O => \N__39524\,
            I => \bfn_17_16_0_\
        );

    \I__8817\ : InMux
    port map (
            O => \N__39521\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__8816\ : CascadeMux
    port map (
            O => \N__39518\,
            I => \N__39515\
        );

    \I__8815\ : InMux
    port map (
            O => \N__39515\,
            I => \N__39512\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__39512\,
            I => \N__39509\
        );

    \I__8813\ : Span4Mux_h
    port map (
            O => \N__39509\,
            I => \N__39506\
        );

    \I__8812\ : Odrv4
    port map (
            O => \N__39506\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__8811\ : InMux
    port map (
            O => \N__39503\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__8810\ : InMux
    port map (
            O => \N__39500\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__8809\ : InMux
    port map (
            O => \N__39497\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__8808\ : InMux
    port map (
            O => \N__39494\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__8807\ : InMux
    port map (
            O => \N__39491\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__8806\ : InMux
    port map (
            O => \N__39488\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__8805\ : InMux
    port map (
            O => \N__39485\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__8804\ : InMux
    port map (
            O => \N__39482\,
            I => \bfn_17_15_0_\
        );

    \I__8803\ : InMux
    port map (
            O => \N__39479\,
            I => \N__39473\
        );

    \I__8802\ : InMux
    port map (
            O => \N__39478\,
            I => \N__39473\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__39473\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__8800\ : InMux
    port map (
            O => \N__39470\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__8799\ : InMux
    port map (
            O => \N__39467\,
            I => \N__39463\
        );

    \I__8798\ : InMux
    port map (
            O => \N__39466\,
            I => \N__39460\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__39463\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__39460\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__8795\ : InMux
    port map (
            O => \N__39455\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__8794\ : InMux
    port map (
            O => \N__39452\,
            I => \N__39448\
        );

    \I__8793\ : InMux
    port map (
            O => \N__39451\,
            I => \N__39445\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__39448\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__39445\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__8790\ : InMux
    port map (
            O => \N__39440\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__8789\ : CascadeMux
    port map (
            O => \N__39437\,
            I => \N__39433\
        );

    \I__8788\ : InMux
    port map (
            O => \N__39436\,
            I => \N__39428\
        );

    \I__8787\ : InMux
    port map (
            O => \N__39433\,
            I => \N__39428\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__39428\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__8785\ : InMux
    port map (
            O => \N__39425\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__8784\ : InMux
    port map (
            O => \N__39422\,
            I => \N__39416\
        );

    \I__8783\ : InMux
    port map (
            O => \N__39421\,
            I => \N__39416\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__39416\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__8781\ : InMux
    port map (
            O => \N__39413\,
            I => \bfn_17_13_0_\
        );

    \I__8780\ : InMux
    port map (
            O => \N__39410\,
            I => \N__39407\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__39407\,
            I => \N__39403\
        );

    \I__8778\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39400\
        );

    \I__8777\ : Odrv4
    port map (
            O => \N__39403\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__39400\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__8775\ : InMux
    port map (
            O => \N__39395\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__8774\ : InMux
    port map (
            O => \N__39392\,
            I => \N__39389\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__39389\,
            I => \N__39385\
        );

    \I__8772\ : CascadeMux
    port map (
            O => \N__39388\,
            I => \N__39382\
        );

    \I__8771\ : Span4Mux_h
    port map (
            O => \N__39385\,
            I => \N__39379\
        );

    \I__8770\ : InMux
    port map (
            O => \N__39382\,
            I => \N__39376\
        );

    \I__8769\ : Odrv4
    port map (
            O => \N__39379\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__39376\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__8767\ : InMux
    port map (
            O => \N__39371\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__8766\ : InMux
    port map (
            O => \N__39368\,
            I => \N__39365\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__39365\,
            I => \N__39362\
        );

    \I__8764\ : Span4Mux_h
    port map (
            O => \N__39362\,
            I => \N__39358\
        );

    \I__8763\ : InMux
    port map (
            O => \N__39361\,
            I => \N__39355\
        );

    \I__8762\ : Odrv4
    port map (
            O => \N__39358\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__39355\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__8760\ : InMux
    port map (
            O => \N__39350\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__8759\ : InMux
    port map (
            O => \N__39347\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__8758\ : InMux
    port map (
            O => \N__39344\,
            I => \N__39339\
        );

    \I__8757\ : InMux
    port map (
            O => \N__39343\,
            I => \N__39334\
        );

    \I__8756\ : InMux
    port map (
            O => \N__39342\,
            I => \N__39331\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__39339\,
            I => \N__39328\
        );

    \I__8754\ : InMux
    port map (
            O => \N__39338\,
            I => \N__39325\
        );

    \I__8753\ : InMux
    port map (
            O => \N__39337\,
            I => \N__39322\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__39334\,
            I => \N__39319\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__39331\,
            I => \N__39316\
        );

    \I__8750\ : Span4Mux_h
    port map (
            O => \N__39328\,
            I => \N__39313\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__39325\,
            I => \N__39308\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__39322\,
            I => \N__39308\
        );

    \I__8747\ : Span4Mux_h
    port map (
            O => \N__39319\,
            I => \N__39303\
        );

    \I__8746\ : Span4Mux_h
    port map (
            O => \N__39316\,
            I => \N__39303\
        );

    \I__8745\ : Odrv4
    port map (
            O => \N__39313\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__8744\ : Odrv12
    port map (
            O => \N__39308\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__8743\ : Odrv4
    port map (
            O => \N__39303\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__8742\ : CEMux
    port map (
            O => \N__39296\,
            I => \N__39278\
        );

    \I__8741\ : CEMux
    port map (
            O => \N__39295\,
            I => \N__39278\
        );

    \I__8740\ : CEMux
    port map (
            O => \N__39294\,
            I => \N__39278\
        );

    \I__8739\ : CEMux
    port map (
            O => \N__39293\,
            I => \N__39278\
        );

    \I__8738\ : CEMux
    port map (
            O => \N__39292\,
            I => \N__39278\
        );

    \I__8737\ : CEMux
    port map (
            O => \N__39291\,
            I => \N__39278\
        );

    \I__8736\ : GlobalMux
    port map (
            O => \N__39278\,
            I => \N__39275\
        );

    \I__8735\ : gio2CtrlBuf
    port map (
            O => \N__39275\,
            I => \delay_measurement_inst.delay_tr_timer.N_434_i_g\
        );

    \I__8734\ : InMux
    port map (
            O => \N__39272\,
            I => \N__39269\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__39269\,
            I => \N__39265\
        );

    \I__8732\ : InMux
    port map (
            O => \N__39268\,
            I => \N__39262\
        );

    \I__8731\ : Span4Mux_v
    port map (
            O => \N__39265\,
            I => \N__39256\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__39262\,
            I => \N__39256\
        );

    \I__8729\ : InMux
    port map (
            O => \N__39261\,
            I => \N__39253\
        );

    \I__8728\ : Odrv4
    port map (
            O => \N__39256\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__39253\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__8726\ : InMux
    port map (
            O => \N__39248\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__8725\ : CascadeMux
    port map (
            O => \N__39245\,
            I => \N__39242\
        );

    \I__8724\ : InMux
    port map (
            O => \N__39242\,
            I => \N__39239\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__39239\,
            I => \N__39235\
        );

    \I__8722\ : CascadeMux
    port map (
            O => \N__39238\,
            I => \N__39231\
        );

    \I__8721\ : Span4Mux_v
    port map (
            O => \N__39235\,
            I => \N__39228\
        );

    \I__8720\ : InMux
    port map (
            O => \N__39234\,
            I => \N__39225\
        );

    \I__8719\ : InMux
    port map (
            O => \N__39231\,
            I => \N__39222\
        );

    \I__8718\ : Odrv4
    port map (
            O => \N__39228\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__39225\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__39222\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__8715\ : InMux
    port map (
            O => \N__39215\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__8714\ : InMux
    port map (
            O => \N__39212\,
            I => \N__39209\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__39209\,
            I => \N__39206\
        );

    \I__8712\ : Span4Mux_v
    port map (
            O => \N__39206\,
            I => \N__39201\
        );

    \I__8711\ : InMux
    port map (
            O => \N__39205\,
            I => \N__39196\
        );

    \I__8710\ : InMux
    port map (
            O => \N__39204\,
            I => \N__39196\
        );

    \I__8709\ : Odrv4
    port map (
            O => \N__39201\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__39196\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__8707\ : InMux
    port map (
            O => \N__39191\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__8706\ : InMux
    port map (
            O => \N__39188\,
            I => \N__39185\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__39185\,
            I => \N__39181\
        );

    \I__8704\ : CascadeMux
    port map (
            O => \N__39184\,
            I => \N__39178\
        );

    \I__8703\ : Span4Mux_v
    port map (
            O => \N__39181\,
            I => \N__39174\
        );

    \I__8702\ : InMux
    port map (
            O => \N__39178\,
            I => \N__39169\
        );

    \I__8701\ : InMux
    port map (
            O => \N__39177\,
            I => \N__39169\
        );

    \I__8700\ : Odrv4
    port map (
            O => \N__39174\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__39169\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__8698\ : InMux
    port map (
            O => \N__39164\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__8697\ : InMux
    port map (
            O => \N__39161\,
            I => \N__39158\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__39158\,
            I => \N__39153\
        );

    \I__8695\ : InMux
    port map (
            O => \N__39157\,
            I => \N__39148\
        );

    \I__8694\ : InMux
    port map (
            O => \N__39156\,
            I => \N__39148\
        );

    \I__8693\ : Span4Mux_v
    port map (
            O => \N__39153\,
            I => \N__39145\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__39148\,
            I => \N__39142\
        );

    \I__8691\ : Odrv4
    port map (
            O => \N__39145\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__8690\ : Odrv4
    port map (
            O => \N__39142\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__8689\ : InMux
    port map (
            O => \N__39137\,
            I => \bfn_17_12_0_\
        );

    \I__8688\ : InMux
    port map (
            O => \N__39134\,
            I => \N__39131\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__39131\,
            I => \N__39127\
        );

    \I__8686\ : InMux
    port map (
            O => \N__39130\,
            I => \N__39124\
        );

    \I__8685\ : Odrv12
    port map (
            O => \N__39127\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__39124\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__8683\ : InMux
    port map (
            O => \N__39119\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__8682\ : CascadeMux
    port map (
            O => \N__39116\,
            I => \N__39113\
        );

    \I__8681\ : InMux
    port map (
            O => \N__39113\,
            I => \N__39109\
        );

    \I__8680\ : InMux
    port map (
            O => \N__39112\,
            I => \N__39106\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__39109\,
            I => \N__39103\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__39106\,
            I => \N__39100\
        );

    \I__8677\ : Odrv12
    port map (
            O => \N__39103\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__8676\ : Odrv4
    port map (
            O => \N__39100\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__8675\ : InMux
    port map (
            O => \N__39095\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__8674\ : InMux
    port map (
            O => \N__39092\,
            I => \N__39088\
        );

    \I__8673\ : CascadeMux
    port map (
            O => \N__39091\,
            I => \N__39085\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__39088\,
            I => \N__39082\
        );

    \I__8671\ : InMux
    port map (
            O => \N__39085\,
            I => \N__39079\
        );

    \I__8670\ : Sp12to4
    port map (
            O => \N__39082\,
            I => \N__39074\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__39079\,
            I => \N__39074\
        );

    \I__8668\ : Odrv12
    port map (
            O => \N__39074\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__8667\ : InMux
    port map (
            O => \N__39071\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__8666\ : InMux
    port map (
            O => \N__39068\,
            I => \N__39065\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__39065\,
            I => \N__39062\
        );

    \I__8664\ : Span4Mux_v
    port map (
            O => \N__39062\,
            I => \N__39057\
        );

    \I__8663\ : InMux
    port map (
            O => \N__39061\,
            I => \N__39052\
        );

    \I__8662\ : InMux
    port map (
            O => \N__39060\,
            I => \N__39052\
        );

    \I__8661\ : Odrv4
    port map (
            O => \N__39057\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__39052\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__8659\ : InMux
    port map (
            O => \N__39047\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__8658\ : CascadeMux
    port map (
            O => \N__39044\,
            I => \N__39041\
        );

    \I__8657\ : InMux
    port map (
            O => \N__39041\,
            I => \N__39038\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__39038\,
            I => \N__39034\
        );

    \I__8655\ : CascadeMux
    port map (
            O => \N__39037\,
            I => \N__39030\
        );

    \I__8654\ : Span4Mux_h
    port map (
            O => \N__39034\,
            I => \N__39027\
        );

    \I__8653\ : InMux
    port map (
            O => \N__39033\,
            I => \N__39024\
        );

    \I__8652\ : InMux
    port map (
            O => \N__39030\,
            I => \N__39021\
        );

    \I__8651\ : Odrv4
    port map (
            O => \N__39027\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__39024\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__39021\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__8648\ : InMux
    port map (
            O => \N__39014\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__8647\ : CascadeMux
    port map (
            O => \N__39011\,
            I => \N__39008\
        );

    \I__8646\ : InMux
    port map (
            O => \N__39008\,
            I => \N__39005\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__39005\,
            I => \N__39001\
        );

    \I__8644\ : CascadeMux
    port map (
            O => \N__39004\,
            I => \N__38996\
        );

    \I__8643\ : Span4Mux_v
    port map (
            O => \N__39001\,
            I => \N__38993\
        );

    \I__8642\ : InMux
    port map (
            O => \N__39000\,
            I => \N__38990\
        );

    \I__8641\ : InMux
    port map (
            O => \N__38999\,
            I => \N__38985\
        );

    \I__8640\ : InMux
    port map (
            O => \N__38996\,
            I => \N__38985\
        );

    \I__8639\ : Odrv4
    port map (
            O => \N__38993\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__38990\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__38985\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__8636\ : InMux
    port map (
            O => \N__38978\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__8635\ : InMux
    port map (
            O => \N__38975\,
            I => \N__38972\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__38972\,
            I => \N__38969\
        );

    \I__8633\ : Span4Mux_h
    port map (
            O => \N__38969\,
            I => \N__38965\
        );

    \I__8632\ : InMux
    port map (
            O => \N__38968\,
            I => \N__38962\
        );

    \I__8631\ : Odrv4
    port map (
            O => \N__38965\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__38962\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__8629\ : InMux
    port map (
            O => \N__38957\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__8628\ : InMux
    port map (
            O => \N__38954\,
            I => \N__38951\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__38951\,
            I => \N__38948\
        );

    \I__8626\ : Span4Mux_h
    port map (
            O => \N__38948\,
            I => \N__38944\
        );

    \I__8625\ : InMux
    port map (
            O => \N__38947\,
            I => \N__38941\
        );

    \I__8624\ : Odrv4
    port map (
            O => \N__38944\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__38941\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__8622\ : InMux
    port map (
            O => \N__38936\,
            I => \bfn_17_11_0_\
        );

    \I__8621\ : InMux
    port map (
            O => \N__38933\,
            I => \N__38930\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__38930\,
            I => \N__38927\
        );

    \I__8619\ : Span4Mux_h
    port map (
            O => \N__38927\,
            I => \N__38923\
        );

    \I__8618\ : InMux
    port map (
            O => \N__38926\,
            I => \N__38920\
        );

    \I__8617\ : Odrv4
    port map (
            O => \N__38923\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__38920\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__8615\ : InMux
    port map (
            O => \N__38915\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__8614\ : InMux
    port map (
            O => \N__38912\,
            I => \N__38909\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__38909\,
            I => \N__38905\
        );

    \I__8612\ : CascadeMux
    port map (
            O => \N__38908\,
            I => \N__38902\
        );

    \I__8611\ : Span4Mux_v
    port map (
            O => \N__38905\,
            I => \N__38899\
        );

    \I__8610\ : InMux
    port map (
            O => \N__38902\,
            I => \N__38896\
        );

    \I__8609\ : Odrv4
    port map (
            O => \N__38899\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__38896\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__8607\ : InMux
    port map (
            O => \N__38891\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__8606\ : CascadeMux
    port map (
            O => \N__38888\,
            I => \N__38884\
        );

    \I__8605\ : CascadeMux
    port map (
            O => \N__38887\,
            I => \N__38881\
        );

    \I__8604\ : InMux
    port map (
            O => \N__38884\,
            I => \N__38878\
        );

    \I__8603\ : InMux
    port map (
            O => \N__38881\,
            I => \N__38875\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__38878\,
            I => \N__38870\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__38875\,
            I => \N__38867\
        );

    \I__8600\ : InMux
    port map (
            O => \N__38874\,
            I => \N__38862\
        );

    \I__8599\ : InMux
    port map (
            O => \N__38873\,
            I => \N__38862\
        );

    \I__8598\ : Odrv4
    port map (
            O => \N__38870\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__8597\ : Odrv4
    port map (
            O => \N__38867\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__38862\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__8595\ : InMux
    port map (
            O => \N__38855\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__8594\ : InMux
    port map (
            O => \N__38852\,
            I => \N__38849\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__38849\,
            I => \N__38846\
        );

    \I__8592\ : Span4Mux_h
    port map (
            O => \N__38846\,
            I => \N__38843\
        );

    \I__8591\ : Odrv4
    port map (
            O => \N__38843\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__8590\ : InMux
    port map (
            O => \N__38840\,
            I => \N__38834\
        );

    \I__8589\ : InMux
    port map (
            O => \N__38839\,
            I => \N__38834\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__38834\,
            I => \N__38831\
        );

    \I__8587\ : Span4Mux_v
    port map (
            O => \N__38831\,
            I => \N__38827\
        );

    \I__8586\ : InMux
    port map (
            O => \N__38830\,
            I => \N__38824\
        );

    \I__8585\ : Odrv4
    port map (
            O => \N__38827\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__38824\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__8583\ : InMux
    port map (
            O => \N__38819\,
            I => \N__38815\
        );

    \I__8582\ : InMux
    port map (
            O => \N__38818\,
            I => \N__38812\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__38815\,
            I => \N__38807\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__38812\,
            I => \N__38807\
        );

    \I__8579\ : Odrv4
    port map (
            O => \N__38807\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__8578\ : InMux
    port map (
            O => \N__38804\,
            I => \N__38801\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__38801\,
            I => \N__38797\
        );

    \I__8576\ : InMux
    port map (
            O => \N__38800\,
            I => \N__38794\
        );

    \I__8575\ : Span4Mux_v
    port map (
            O => \N__38797\,
            I => \N__38788\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__38794\,
            I => \N__38788\
        );

    \I__8573\ : InMux
    port map (
            O => \N__38793\,
            I => \N__38785\
        );

    \I__8572\ : Span4Mux_v
    port map (
            O => \N__38788\,
            I => \N__38780\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__38785\,
            I => \N__38780\
        );

    \I__8570\ : Span4Mux_h
    port map (
            O => \N__38780\,
            I => \N__38777\
        );

    \I__8569\ : Odrv4
    port map (
            O => \N__38777\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__8568\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38771\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__38771\,
            I => \N__38767\
        );

    \I__8566\ : InMux
    port map (
            O => \N__38770\,
            I => \N__38764\
        );

    \I__8565\ : Odrv4
    port map (
            O => \N__38767\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__38764\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__8563\ : InMux
    port map (
            O => \N__38759\,
            I => \N__38756\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__38756\,
            I => \N__38753\
        );

    \I__8561\ : Span4Mux_h
    port map (
            O => \N__38753\,
            I => \N__38750\
        );

    \I__8560\ : Odrv4
    port map (
            O => \N__38750\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__8559\ : InMux
    port map (
            O => \N__38747\,
            I => \N__38743\
        );

    \I__8558\ : InMux
    port map (
            O => \N__38746\,
            I => \N__38740\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__38743\,
            I => \N__38736\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__38740\,
            I => \N__38733\
        );

    \I__8555\ : InMux
    port map (
            O => \N__38739\,
            I => \N__38730\
        );

    \I__8554\ : Span4Mux_v
    port map (
            O => \N__38736\,
            I => \N__38727\
        );

    \I__8553\ : Span4Mux_h
    port map (
            O => \N__38733\,
            I => \N__38722\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__38730\,
            I => \N__38722\
        );

    \I__8551\ : Odrv4
    port map (
            O => \N__38727\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__8550\ : Odrv4
    port map (
            O => \N__38722\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__8549\ : InMux
    port map (
            O => \N__38717\,
            I => \N__38714\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__38714\,
            I => \N__38711\
        );

    \I__8547\ : Span4Mux_v
    port map (
            O => \N__38711\,
            I => \N__38707\
        );

    \I__8546\ : InMux
    port map (
            O => \N__38710\,
            I => \N__38704\
        );

    \I__8545\ : Odrv4
    port map (
            O => \N__38707\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__38704\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__8543\ : CascadeMux
    port map (
            O => \N__38699\,
            I => \N__38696\
        );

    \I__8542\ : InMux
    port map (
            O => \N__38696\,
            I => \N__38693\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__38693\,
            I => \N__38690\
        );

    \I__8540\ : Span4Mux_v
    port map (
            O => \N__38690\,
            I => \N__38687\
        );

    \I__8539\ : Odrv4
    port map (
            O => \N__38687\,
            I => \current_shift_inst.un38_control_input_cry_18_c_RNOZ0\
        );

    \I__8538\ : CascadeMux
    port map (
            O => \N__38684\,
            I => \N__38681\
        );

    \I__8537\ : InMux
    port map (
            O => \N__38681\,
            I => \N__38678\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__38678\,
            I => \N__38675\
        );

    \I__8535\ : Span4Mux_h
    port map (
            O => \N__38675\,
            I => \N__38672\
        );

    \I__8534\ : Span4Mux_v
    port map (
            O => \N__38672\,
            I => \N__38668\
        );

    \I__8533\ : InMux
    port map (
            O => \N__38671\,
            I => \N__38665\
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__38668\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__38665\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__8530\ : CascadeMux
    port map (
            O => \N__38660\,
            I => \N__38657\
        );

    \I__8529\ : InMux
    port map (
            O => \N__38657\,
            I => \N__38654\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__38654\,
            I => \N__38651\
        );

    \I__8527\ : Span4Mux_v
    port map (
            O => \N__38651\,
            I => \N__38647\
        );

    \I__8526\ : CascadeMux
    port map (
            O => \N__38650\,
            I => \N__38643\
        );

    \I__8525\ : Span4Mux_h
    port map (
            O => \N__38647\,
            I => \N__38640\
        );

    \I__8524\ : InMux
    port map (
            O => \N__38646\,
            I => \N__38637\
        );

    \I__8523\ : InMux
    port map (
            O => \N__38643\,
            I => \N__38634\
        );

    \I__8522\ : Odrv4
    port map (
            O => \N__38640\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__38637\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__38634\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__8519\ : InMux
    port map (
            O => \N__38627\,
            I => \N__38624\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__38624\,
            I => \N__38621\
        );

    \I__8517\ : Span4Mux_v
    port map (
            O => \N__38621\,
            I => \N__38617\
        );

    \I__8516\ : InMux
    port map (
            O => \N__38620\,
            I => \N__38614\
        );

    \I__8515\ : Odrv4
    port map (
            O => \N__38617\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__38614\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__8513\ : InMux
    port map (
            O => \N__38609\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__8512\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38603\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__38603\,
            I => \N__38600\
        );

    \I__8510\ : Span4Mux_h
    port map (
            O => \N__38600\,
            I => \N__38597\
        );

    \I__8509\ : Span4Mux_v
    port map (
            O => \N__38597\,
            I => \N__38593\
        );

    \I__8508\ : InMux
    port map (
            O => \N__38596\,
            I => \N__38590\
        );

    \I__8507\ : Odrv4
    port map (
            O => \N__38593\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__38590\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__8505\ : InMux
    port map (
            O => \N__38585\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__8504\ : CascadeMux
    port map (
            O => \N__38582\,
            I => \N__38579\
        );

    \I__8503\ : InMux
    port map (
            O => \N__38579\,
            I => \N__38576\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__38576\,
            I => \N__38573\
        );

    \I__8501\ : Span4Mux_v
    port map (
            O => \N__38573\,
            I => \N__38567\
        );

    \I__8500\ : InMux
    port map (
            O => \N__38572\,
            I => \N__38562\
        );

    \I__8499\ : InMux
    port map (
            O => \N__38571\,
            I => \N__38562\
        );

    \I__8498\ : InMux
    port map (
            O => \N__38570\,
            I => \N__38559\
        );

    \I__8497\ : Odrv4
    port map (
            O => \N__38567\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__38562\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__38559\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__8494\ : InMux
    port map (
            O => \N__38552\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__8493\ : InMux
    port map (
            O => \N__38549\,
            I => \N__38545\
        );

    \I__8492\ : InMux
    port map (
            O => \N__38548\,
            I => \N__38542\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__38545\,
            I => \N__38537\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__38542\,
            I => \N__38537\
        );

    \I__8489\ : Span4Mux_v
    port map (
            O => \N__38537\,
            I => \N__38533\
        );

    \I__8488\ : InMux
    port map (
            O => \N__38536\,
            I => \N__38530\
        );

    \I__8487\ : Odrv4
    port map (
            O => \N__38533\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__38530\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__8485\ : InMux
    port map (
            O => \N__38525\,
            I => \N__38521\
        );

    \I__8484\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38518\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__38521\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__38518\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__8481\ : InMux
    port map (
            O => \N__38513\,
            I => \N__38509\
        );

    \I__8480\ : InMux
    port map (
            O => \N__38512\,
            I => \N__38505\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__38509\,
            I => \N__38502\
        );

    \I__8478\ : InMux
    port map (
            O => \N__38508\,
            I => \N__38499\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__38505\,
            I => \N__38492\
        );

    \I__8476\ : Span4Mux_v
    port map (
            O => \N__38502\,
            I => \N__38492\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__38499\,
            I => \N__38492\
        );

    \I__8474\ : Odrv4
    port map (
            O => \N__38492\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__8473\ : InMux
    port map (
            O => \N__38489\,
            I => \N__38485\
        );

    \I__8472\ : InMux
    port map (
            O => \N__38488\,
            I => \N__38482\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__38485\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__38482\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__8469\ : InMux
    port map (
            O => \N__38477\,
            I => \N__38474\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__38474\,
            I => \N__38469\
        );

    \I__8467\ : InMux
    port map (
            O => \N__38473\,
            I => \N__38464\
        );

    \I__8466\ : InMux
    port map (
            O => \N__38472\,
            I => \N__38464\
        );

    \I__8465\ : Odrv12
    port map (
            O => \N__38469\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__38464\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__8463\ : InMux
    port map (
            O => \N__38459\,
            I => \N__38456\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__38456\,
            I => \N__38452\
        );

    \I__8461\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38449\
        );

    \I__8460\ : Odrv4
    port map (
            O => \N__38452\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__38449\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__8458\ : InMux
    port map (
            O => \N__38444\,
            I => \N__38441\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__38441\,
            I => \N__38438\
        );

    \I__8456\ : Odrv12
    port map (
            O => \N__38438\,
            I => \current_shift_inst.un38_control_input_cry_16_c_RNOZ0\
        );

    \I__8455\ : InMux
    port map (
            O => \N__38435\,
            I => \N__38432\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__38432\,
            I => \N__38428\
        );

    \I__8453\ : InMux
    port map (
            O => \N__38431\,
            I => \N__38425\
        );

    \I__8452\ : Span4Mux_v
    port map (
            O => \N__38428\,
            I => \N__38422\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__38425\,
            I => \N__38419\
        );

    \I__8450\ : Span4Mux_v
    port map (
            O => \N__38422\,
            I => \N__38415\
        );

    \I__8449\ : Span4Mux_h
    port map (
            O => \N__38419\,
            I => \N__38412\
        );

    \I__8448\ : InMux
    port map (
            O => \N__38418\,
            I => \N__38409\
        );

    \I__8447\ : Odrv4
    port map (
            O => \N__38415\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8446\ : Odrv4
    port map (
            O => \N__38412\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__38409\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__8444\ : InMux
    port map (
            O => \N__38402\,
            I => \N__38399\
        );

    \I__8443\ : LocalMux
    port map (
            O => \N__38399\,
            I => \N__38396\
        );

    \I__8442\ : Span4Mux_h
    port map (
            O => \N__38396\,
            I => \N__38392\
        );

    \I__8441\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38389\
        );

    \I__8440\ : Odrv4
    port map (
            O => \N__38392\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__38389\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8438\ : InMux
    port map (
            O => \N__38384\,
            I => \N__38380\
        );

    \I__8437\ : InMux
    port map (
            O => \N__38383\,
            I => \N__38377\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__38380\,
            I => \N__38374\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__38377\,
            I => \N__38370\
        );

    \I__8434\ : Span4Mux_h
    port map (
            O => \N__38374\,
            I => \N__38367\
        );

    \I__8433\ : InMux
    port map (
            O => \N__38373\,
            I => \N__38364\
        );

    \I__8432\ : Odrv12
    port map (
            O => \N__38370\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8431\ : Odrv4
    port map (
            O => \N__38367\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__38364\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__8429\ : InMux
    port map (
            O => \N__38357\,
            I => \N__38354\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__38354\,
            I => \N__38350\
        );

    \I__8427\ : InMux
    port map (
            O => \N__38353\,
            I => \N__38347\
        );

    \I__8426\ : Odrv4
    port map (
            O => \N__38350\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__38347\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8424\ : InMux
    port map (
            O => \N__38342\,
            I => \N__38339\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__38339\,
            I => \N__38336\
        );

    \I__8422\ : Span4Mux_h
    port map (
            O => \N__38336\,
            I => \N__38333\
        );

    \I__8421\ : Span4Mux_h
    port map (
            O => \N__38333\,
            I => \N__38330\
        );

    \I__8420\ : Odrv4
    port map (
            O => \N__38330\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__8419\ : InMux
    port map (
            O => \N__38327\,
            I => \N__38324\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__38324\,
            I => \N__38321\
        );

    \I__8417\ : Span4Mux_h
    port map (
            O => \N__38321\,
            I => \N__38318\
        );

    \I__8416\ : Span4Mux_v
    port map (
            O => \N__38318\,
            I => \N__38315\
        );

    \I__8415\ : Span4Mux_v
    port map (
            O => \N__38315\,
            I => \N__38312\
        );

    \I__8414\ : Odrv4
    port map (
            O => \N__38312\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__8413\ : InMux
    port map (
            O => \N__38309\,
            I => \N__38305\
        );

    \I__8412\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38302\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__38305\,
            I => \N__38299\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__38302\,
            I => \N__38296\
        );

    \I__8409\ : Span4Mux_v
    port map (
            O => \N__38299\,
            I => \N__38292\
        );

    \I__8408\ : Span4Mux_h
    port map (
            O => \N__38296\,
            I => \N__38289\
        );

    \I__8407\ : InMux
    port map (
            O => \N__38295\,
            I => \N__38286\
        );

    \I__8406\ : Odrv4
    port map (
            O => \N__38292\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8405\ : Odrv4
    port map (
            O => \N__38289\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__38286\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__8403\ : InMux
    port map (
            O => \N__38279\,
            I => \N__38275\
        );

    \I__8402\ : InMux
    port map (
            O => \N__38278\,
            I => \N__38272\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__38275\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__38272\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8399\ : InMux
    port map (
            O => \N__38267\,
            I => \N__38264\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__38264\,
            I => \N__38260\
        );

    \I__8397\ : InMux
    port map (
            O => \N__38263\,
            I => \N__38256\
        );

    \I__8396\ : Span4Mux_v
    port map (
            O => \N__38260\,
            I => \N__38253\
        );

    \I__8395\ : InMux
    port map (
            O => \N__38259\,
            I => \N__38250\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__38256\,
            I => \N__38247\
        );

    \I__8393\ : Sp12to4
    port map (
            O => \N__38253\,
            I => \N__38242\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__38250\,
            I => \N__38242\
        );

    \I__8391\ : Odrv4
    port map (
            O => \N__38247\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__8390\ : Odrv12
    port map (
            O => \N__38242\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__8389\ : InMux
    port map (
            O => \N__38237\,
            I => \N__38233\
        );

    \I__8388\ : InMux
    port map (
            O => \N__38236\,
            I => \N__38230\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__38233\,
            I => \N__38227\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__38230\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__8385\ : Odrv4
    port map (
            O => \N__38227\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__8384\ : InMux
    port map (
            O => \N__38222\,
            I => \N__38219\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__38219\,
            I => \N__38216\
        );

    \I__8382\ : Span4Mux_h
    port map (
            O => \N__38216\,
            I => \N__38213\
        );

    \I__8381\ : Odrv4
    port map (
            O => \N__38213\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__8380\ : InMux
    port map (
            O => \N__38210\,
            I => \N__38204\
        );

    \I__8379\ : InMux
    port map (
            O => \N__38209\,
            I => \N__38204\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__38204\,
            I => \N__38200\
        );

    \I__8377\ : InMux
    port map (
            O => \N__38203\,
            I => \N__38197\
        );

    \I__8376\ : Span4Mux_h
    port map (
            O => \N__38200\,
            I => \N__38194\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__38197\,
            I => \N__38191\
        );

    \I__8374\ : Span4Mux_v
    port map (
            O => \N__38194\,
            I => \N__38188\
        );

    \I__8373\ : Span4Mux_v
    port map (
            O => \N__38191\,
            I => \N__38185\
        );

    \I__8372\ : Odrv4
    port map (
            O => \N__38188\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__8371\ : Odrv4
    port map (
            O => \N__38185\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__8370\ : CEMux
    port map (
            O => \N__38180\,
            I => \N__38162\
        );

    \I__8369\ : CEMux
    port map (
            O => \N__38179\,
            I => \N__38162\
        );

    \I__8368\ : CEMux
    port map (
            O => \N__38178\,
            I => \N__38162\
        );

    \I__8367\ : CEMux
    port map (
            O => \N__38177\,
            I => \N__38162\
        );

    \I__8366\ : CEMux
    port map (
            O => \N__38176\,
            I => \N__38162\
        );

    \I__8365\ : CEMux
    port map (
            O => \N__38175\,
            I => \N__38162\
        );

    \I__8364\ : GlobalMux
    port map (
            O => \N__38162\,
            I => \N__38159\
        );

    \I__8363\ : gio2CtrlBuf
    port map (
            O => \N__38159\,
            I => \current_shift_inst.timer_s1.N_166_i_g\
        );

    \I__8362\ : InMux
    port map (
            O => \N__38156\,
            I => \N__38150\
        );

    \I__8361\ : InMux
    port map (
            O => \N__38155\,
            I => \N__38150\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__38150\,
            I => \N__38147\
        );

    \I__8359\ : Span4Mux_v
    port map (
            O => \N__38147\,
            I => \N__38144\
        );

    \I__8358\ : Span4Mux_h
    port map (
            O => \N__38144\,
            I => \N__38140\
        );

    \I__8357\ : InMux
    port map (
            O => \N__38143\,
            I => \N__38137\
        );

    \I__8356\ : Odrv4
    port map (
            O => \N__38140\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__38137\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__8354\ : InMux
    port map (
            O => \N__38132\,
            I => \N__38126\
        );

    \I__8353\ : InMux
    port map (
            O => \N__38131\,
            I => \N__38126\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__38126\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__8351\ : CascadeMux
    port map (
            O => \N__38123\,
            I => \N__38119\
        );

    \I__8350\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38115\
        );

    \I__8349\ : InMux
    port map (
            O => \N__38119\,
            I => \N__38110\
        );

    \I__8348\ : InMux
    port map (
            O => \N__38118\,
            I => \N__38110\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__38115\,
            I => \N__38107\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__38110\,
            I => \N__38104\
        );

    \I__8345\ : Span4Mux_h
    port map (
            O => \N__38107\,
            I => \N__38101\
        );

    \I__8344\ : Span4Mux_h
    port map (
            O => \N__38104\,
            I => \N__38098\
        );

    \I__8343\ : Odrv4
    port map (
            O => \N__38101\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__8342\ : Odrv4
    port map (
            O => \N__38098\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__8341\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38090\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__38090\,
            I => \N__38087\
        );

    \I__8339\ : Span4Mux_v
    port map (
            O => \N__38087\,
            I => \N__38083\
        );

    \I__8338\ : InMux
    port map (
            O => \N__38086\,
            I => \N__38080\
        );

    \I__8337\ : Odrv4
    port map (
            O => \N__38083\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__38080\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__8335\ : InMux
    port map (
            O => \N__38075\,
            I => \N__38069\
        );

    \I__8334\ : InMux
    port map (
            O => \N__38074\,
            I => \N__38069\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__38069\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__8332\ : InMux
    port map (
            O => \N__38066\,
            I => \N__38060\
        );

    \I__8331\ : InMux
    port map (
            O => \N__38065\,
            I => \N__38060\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__38060\,
            I => \N__38057\
        );

    \I__8329\ : Span4Mux_h
    port map (
            O => \N__38057\,
            I => \N__38053\
        );

    \I__8328\ : InMux
    port map (
            O => \N__38056\,
            I => \N__38050\
        );

    \I__8327\ : Odrv4
    port map (
            O => \N__38053\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__38050\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__8325\ : InMux
    port map (
            O => \N__38045\,
            I => \N__38042\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__38042\,
            I => \N__38039\
        );

    \I__8323\ : Span4Mux_h
    port map (
            O => \N__38039\,
            I => \N__38036\
        );

    \I__8322\ : Odrv4
    port map (
            O => \N__38036\,
            I => \current_shift_inst.un38_control_input_cry_17_c_RNOZ0\
        );

    \I__8321\ : InMux
    port map (
            O => \N__38033\,
            I => \N__38030\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__38030\,
            I => \N__38026\
        );

    \I__8319\ : InMux
    port map (
            O => \N__38029\,
            I => \N__38023\
        );

    \I__8318\ : Span4Mux_v
    port map (
            O => \N__38026\,
            I => \N__38018\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__38023\,
            I => \N__38018\
        );

    \I__8316\ : Span4Mux_h
    port map (
            O => \N__38018\,
            I => \N__38014\
        );

    \I__8315\ : InMux
    port map (
            O => \N__38017\,
            I => \N__38011\
        );

    \I__8314\ : Odrv4
    port map (
            O => \N__38014\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__38011\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__8312\ : InMux
    port map (
            O => \N__38006\,
            I => \N__38003\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__38003\,
            I => \N__37999\
        );

    \I__8310\ : InMux
    port map (
            O => \N__38002\,
            I => \N__37996\
        );

    \I__8309\ : Odrv4
    port map (
            O => \N__37999\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__37996\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__8307\ : CascadeMux
    port map (
            O => \N__37991\,
            I => \N__37988\
        );

    \I__8306\ : InMux
    port map (
            O => \N__37988\,
            I => \N__37985\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__37985\,
            I => \N__37982\
        );

    \I__8304\ : Span12Mux_v
    port map (
            O => \N__37982\,
            I => \N__37979\
        );

    \I__8303\ : Odrv12
    port map (
            O => \N__37979\,
            I => \current_shift_inst.un38_control_input_cry_14_c_RNOZ0\
        );

    \I__8302\ : InMux
    port map (
            O => \N__37976\,
            I => \N__37972\
        );

    \I__8301\ : InMux
    port map (
            O => \N__37975\,
            I => \N__37969\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__37972\,
            I => \N__37966\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__37969\,
            I => \N__37963\
        );

    \I__8298\ : Span4Mux_h
    port map (
            O => \N__37966\,
            I => \N__37957\
        );

    \I__8297\ : Span4Mux_h
    port map (
            O => \N__37963\,
            I => \N__37957\
        );

    \I__8296\ : InMux
    port map (
            O => \N__37962\,
            I => \N__37954\
        );

    \I__8295\ : Odrv4
    port map (
            O => \N__37957\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__37954\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8293\ : InMux
    port map (
            O => \N__37949\,
            I => \N__37946\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__37946\,
            I => \N__37942\
        );

    \I__8291\ : InMux
    port map (
            O => \N__37945\,
            I => \N__37939\
        );

    \I__8290\ : Odrv4
    port map (
            O => \N__37942\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__37939\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8288\ : InMux
    port map (
            O => \N__37934\,
            I => \N__37930\
        );

    \I__8287\ : InMux
    port map (
            O => \N__37933\,
            I => \N__37927\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__37930\,
            I => \N__37924\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__37927\,
            I => \N__37921\
        );

    \I__8284\ : Span4Mux_h
    port map (
            O => \N__37924\,
            I => \N__37917\
        );

    \I__8283\ : Span4Mux_h
    port map (
            O => \N__37921\,
            I => \N__37914\
        );

    \I__8282\ : InMux
    port map (
            O => \N__37920\,
            I => \N__37911\
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__37917\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__8280\ : Odrv4
    port map (
            O => \N__37914\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__37911\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__8278\ : InMux
    port map (
            O => \N__37904\,
            I => \N__37900\
        );

    \I__8277\ : InMux
    port map (
            O => \N__37903\,
            I => \N__37897\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__37900\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__37897\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__8274\ : InMux
    port map (
            O => \N__37892\,
            I => \N__37888\
        );

    \I__8273\ : InMux
    port map (
            O => \N__37891\,
            I => \N__37885\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__37888\,
            I => \N__37882\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__37885\,
            I => \N__37878\
        );

    \I__8270\ : Span4Mux_v
    port map (
            O => \N__37882\,
            I => \N__37875\
        );

    \I__8269\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37872\
        );

    \I__8268\ : Odrv4
    port map (
            O => \N__37878\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__8267\ : Odrv4
    port map (
            O => \N__37875\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__37872\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__8265\ : InMux
    port map (
            O => \N__37865\,
            I => \N__37861\
        );

    \I__8264\ : InMux
    port map (
            O => \N__37864\,
            I => \N__37858\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__37861\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__37858\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__8261\ : InMux
    port map (
            O => \N__37853\,
            I => \N__37850\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__37850\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__8259\ : InMux
    port map (
            O => \N__37847\,
            I => \N__37843\
        );

    \I__8258\ : InMux
    port map (
            O => \N__37846\,
            I => \N__37840\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__37843\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__37840\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__8255\ : InMux
    port map (
            O => \N__37835\,
            I => \N__37830\
        );

    \I__8254\ : InMux
    port map (
            O => \N__37834\,
            I => \N__37825\
        );

    \I__8253\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37825\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__37830\,
            I => \N__37822\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__37825\,
            I => \N__37819\
        );

    \I__8250\ : Span4Mux_v
    port map (
            O => \N__37822\,
            I => \N__37816\
        );

    \I__8249\ : Span4Mux_h
    port map (
            O => \N__37819\,
            I => \N__37813\
        );

    \I__8248\ : Odrv4
    port map (
            O => \N__37816\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__8247\ : Odrv4
    port map (
            O => \N__37813\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__8246\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37804\
        );

    \I__8245\ : InMux
    port map (
            O => \N__37807\,
            I => \N__37801\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__37804\,
            I => \N__37798\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__37801\,
            I => \N__37795\
        );

    \I__8242\ : Span4Mux_h
    port map (
            O => \N__37798\,
            I => \N__37791\
        );

    \I__8241\ : Span4Mux_h
    port map (
            O => \N__37795\,
            I => \N__37788\
        );

    \I__8240\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37785\
        );

    \I__8239\ : Odrv4
    port map (
            O => \N__37791\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__8238\ : Odrv4
    port map (
            O => \N__37788\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__37785\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__8236\ : InMux
    port map (
            O => \N__37778\,
            I => \N__37774\
        );

    \I__8235\ : InMux
    port map (
            O => \N__37777\,
            I => \N__37771\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__37774\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__37771\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__8232\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37763\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__37763\,
            I => \N__37759\
        );

    \I__8230\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37755\
        );

    \I__8229\ : Span4Mux_v
    port map (
            O => \N__37759\,
            I => \N__37752\
        );

    \I__8228\ : InMux
    port map (
            O => \N__37758\,
            I => \N__37749\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__37755\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__8226\ : Odrv4
    port map (
            O => \N__37752\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__37749\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__8224\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37738\
        );

    \I__8223\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37735\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__37738\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__37735\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__8220\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37727\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__37727\,
            I => \N__37717\
        );

    \I__8218\ : InMux
    port map (
            O => \N__37726\,
            I => \N__37702\
        );

    \I__8217\ : InMux
    port map (
            O => \N__37725\,
            I => \N__37702\
        );

    \I__8216\ : InMux
    port map (
            O => \N__37724\,
            I => \N__37702\
        );

    \I__8215\ : InMux
    port map (
            O => \N__37723\,
            I => \N__37702\
        );

    \I__8214\ : InMux
    port map (
            O => \N__37722\,
            I => \N__37702\
        );

    \I__8213\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37702\
        );

    \I__8212\ : InMux
    port map (
            O => \N__37720\,
            I => \N__37702\
        );

    \I__8211\ : Span4Mux_h
    port map (
            O => \N__37717\,
            I => \N__37688\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__37702\,
            I => \N__37688\
        );

    \I__8209\ : InMux
    port map (
            O => \N__37701\,
            I => \N__37673\
        );

    \I__8208\ : InMux
    port map (
            O => \N__37700\,
            I => \N__37673\
        );

    \I__8207\ : InMux
    port map (
            O => \N__37699\,
            I => \N__37673\
        );

    \I__8206\ : InMux
    port map (
            O => \N__37698\,
            I => \N__37673\
        );

    \I__8205\ : InMux
    port map (
            O => \N__37697\,
            I => \N__37673\
        );

    \I__8204\ : InMux
    port map (
            O => \N__37696\,
            I => \N__37673\
        );

    \I__8203\ : InMux
    port map (
            O => \N__37695\,
            I => \N__37673\
        );

    \I__8202\ : InMux
    port map (
            O => \N__37694\,
            I => \N__37668\
        );

    \I__8201\ : InMux
    port map (
            O => \N__37693\,
            I => \N__37668\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__37688\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__37673\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__37668\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8197\ : InMux
    port map (
            O => \N__37661\,
            I => \N__37657\
        );

    \I__8196\ : InMux
    port map (
            O => \N__37660\,
            I => \N__37654\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__37657\,
            I => \N__37651\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__37654\,
            I => \N__37647\
        );

    \I__8193\ : Span4Mux_h
    port map (
            O => \N__37651\,
            I => \N__37644\
        );

    \I__8192\ : InMux
    port map (
            O => \N__37650\,
            I => \N__37641\
        );

    \I__8191\ : Odrv4
    port map (
            O => \N__37647\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__8190\ : Odrv4
    port map (
            O => \N__37644\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__37641\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__8188\ : InMux
    port map (
            O => \N__37634\,
            I => \N__37630\
        );

    \I__8187\ : InMux
    port map (
            O => \N__37633\,
            I => \N__37627\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__37630\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__37627\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__8184\ : InMux
    port map (
            O => \N__37622\,
            I => \N__37609\
        );

    \I__8183\ : InMux
    port map (
            O => \N__37621\,
            I => \N__37609\
        );

    \I__8182\ : InMux
    port map (
            O => \N__37620\,
            I => \N__37609\
        );

    \I__8181\ : InMux
    port map (
            O => \N__37619\,
            I => \N__37606\
        );

    \I__8180\ : InMux
    port map (
            O => \N__37618\,
            I => \N__37599\
        );

    \I__8179\ : InMux
    port map (
            O => \N__37617\,
            I => \N__37599\
        );

    \I__8178\ : InMux
    port map (
            O => \N__37616\,
            I => \N__37599\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__37609\,
            I => \N__37596\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__37606\,
            I => \N__37593\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__37599\,
            I => \N__37582\
        );

    \I__8174\ : Span12Mux_v
    port map (
            O => \N__37596\,
            I => \N__37579\
        );

    \I__8173\ : Span4Mux_h
    port map (
            O => \N__37593\,
            I => \N__37576\
        );

    \I__8172\ : InMux
    port map (
            O => \N__37592\,
            I => \N__37573\
        );

    \I__8171\ : InMux
    port map (
            O => \N__37591\,
            I => \N__37562\
        );

    \I__8170\ : InMux
    port map (
            O => \N__37590\,
            I => \N__37562\
        );

    \I__8169\ : InMux
    port map (
            O => \N__37589\,
            I => \N__37562\
        );

    \I__8168\ : InMux
    port map (
            O => \N__37588\,
            I => \N__37562\
        );

    \I__8167\ : InMux
    port map (
            O => \N__37587\,
            I => \N__37562\
        );

    \I__8166\ : InMux
    port map (
            O => \N__37586\,
            I => \N__37557\
        );

    \I__8165\ : InMux
    port map (
            O => \N__37585\,
            I => \N__37557\
        );

    \I__8164\ : Odrv4
    port map (
            O => \N__37582\,
            I => \phase_controller_inst1.stoper_tr.N_249\
        );

    \I__8163\ : Odrv12
    port map (
            O => \N__37579\,
            I => \phase_controller_inst1.stoper_tr.N_249\
        );

    \I__8162\ : Odrv4
    port map (
            O => \N__37576\,
            I => \phase_controller_inst1.stoper_tr.N_249\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__37573\,
            I => \phase_controller_inst1.stoper_tr.N_249\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__37562\,
            I => \phase_controller_inst1.stoper_tr.N_249\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__37557\,
            I => \phase_controller_inst1.stoper_tr.N_249\
        );

    \I__8158\ : CascadeMux
    port map (
            O => \N__37544\,
            I => \N__37541\
        );

    \I__8157\ : InMux
    port map (
            O => \N__37541\,
            I => \N__37536\
        );

    \I__8156\ : InMux
    port map (
            O => \N__37540\,
            I => \N__37533\
        );

    \I__8155\ : CascadeMux
    port map (
            O => \N__37539\,
            I => \N__37530\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__37536\,
            I => \N__37527\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__37533\,
            I => \N__37524\
        );

    \I__8152\ : InMux
    port map (
            O => \N__37530\,
            I => \N__37520\
        );

    \I__8151\ : Span4Mux_h
    port map (
            O => \N__37527\,
            I => \N__37517\
        );

    \I__8150\ : Sp12to4
    port map (
            O => \N__37524\,
            I => \N__37514\
        );

    \I__8149\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37511\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__37520\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__8147\ : Odrv4
    port map (
            O => \N__37517\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__8146\ : Odrv12
    port map (
            O => \N__37514\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__37511\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__8144\ : CascadeMux
    port map (
            O => \N__37502\,
            I => \N__37499\
        );

    \I__8143\ : InMux
    port map (
            O => \N__37499\,
            I => \N__37494\
        );

    \I__8142\ : CascadeMux
    port map (
            O => \N__37498\,
            I => \N__37489\
        );

    \I__8141\ : CascadeMux
    port map (
            O => \N__37497\,
            I => \N__37485\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__37494\,
            I => \N__37482\
        );

    \I__8139\ : InMux
    port map (
            O => \N__37493\,
            I => \N__37479\
        );

    \I__8138\ : InMux
    port map (
            O => \N__37492\,
            I => \N__37474\
        );

    \I__8137\ : InMux
    port map (
            O => \N__37489\,
            I => \N__37474\
        );

    \I__8136\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37469\
        );

    \I__8135\ : InMux
    port map (
            O => \N__37485\,
            I => \N__37469\
        );

    \I__8134\ : Span4Mux_v
    port map (
            O => \N__37482\,
            I => \N__37466\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__37479\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__37474\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__37469\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2\
        );

    \I__8130\ : Odrv4
    port map (
            O => \N__37466\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2\
        );

    \I__8129\ : InMux
    port map (
            O => \N__37457\,
            I => \N__37454\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__37454\,
            I => \N__37451\
        );

    \I__8127\ : Span4Mux_v
    port map (
            O => \N__37451\,
            I => \N__37446\
        );

    \I__8126\ : InMux
    port map (
            O => \N__37450\,
            I => \N__37441\
        );

    \I__8125\ : InMux
    port map (
            O => \N__37449\,
            I => \N__37441\
        );

    \I__8124\ : Odrv4
    port map (
            O => \N__37446\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__37441\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__8122\ : InMux
    port map (
            O => \N__37436\,
            I => \N__37432\
        );

    \I__8121\ : InMux
    port map (
            O => \N__37435\,
            I => \N__37429\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__37432\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__37429\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__8118\ : InMux
    port map (
            O => \N__37424\,
            I => \N__37421\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__37421\,
            I => \N__37418\
        );

    \I__8116\ : Span4Mux_h
    port map (
            O => \N__37418\,
            I => \N__37415\
        );

    \I__8115\ : Odrv4
    port map (
            O => \N__37415\,
            I => \current_shift_inst.un38_control_input_cry_11_c_RNOZ0\
        );

    \I__8114\ : InMux
    port map (
            O => \N__37412\,
            I => \N__37408\
        );

    \I__8113\ : InMux
    port map (
            O => \N__37411\,
            I => \N__37405\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__37408\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__37405\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8110\ : InMux
    port map (
            O => \N__37400\,
            I => \N__37396\
        );

    \I__8109\ : InMux
    port map (
            O => \N__37399\,
            I => \N__37393\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__37396\,
            I => \N__37388\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__37393\,
            I => \N__37388\
        );

    \I__8106\ : Span4Mux_h
    port map (
            O => \N__37388\,
            I => \N__37384\
        );

    \I__8105\ : InMux
    port map (
            O => \N__37387\,
            I => \N__37381\
        );

    \I__8104\ : Odrv4
    port map (
            O => \N__37384\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__37381\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__8102\ : InMux
    port map (
            O => \N__37376\,
            I => \N__37372\
        );

    \I__8101\ : InMux
    port map (
            O => \N__37375\,
            I => \N__37369\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__37372\,
            I => \N__37364\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__37369\,
            I => \N__37364\
        );

    \I__8098\ : Span4Mux_h
    port map (
            O => \N__37364\,
            I => \N__37360\
        );

    \I__8097\ : InMux
    port map (
            O => \N__37363\,
            I => \N__37357\
        );

    \I__8096\ : Odrv4
    port map (
            O => \N__37360\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__37357\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__8094\ : InMux
    port map (
            O => \N__37352\,
            I => \N__37348\
        );

    \I__8093\ : InMux
    port map (
            O => \N__37351\,
            I => \N__37345\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__37348\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__37345\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8090\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37336\
        );

    \I__8089\ : CascadeMux
    port map (
            O => \N__37339\,
            I => \N__37333\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__37336\,
            I => \N__37329\
        );

    \I__8087\ : InMux
    port map (
            O => \N__37333\,
            I => \N__37324\
        );

    \I__8086\ : InMux
    port map (
            O => \N__37332\,
            I => \N__37324\
        );

    \I__8085\ : Span4Mux_h
    port map (
            O => \N__37329\,
            I => \N__37321\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__37324\,
            I => \N__37318\
        );

    \I__8083\ : Odrv4
    port map (
            O => \N__37321\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__8082\ : Odrv4
    port map (
            O => \N__37318\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__8081\ : InMux
    port map (
            O => \N__37313\,
            I => \N__37309\
        );

    \I__8080\ : InMux
    port map (
            O => \N__37312\,
            I => \N__37306\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__37309\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__37306\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__8077\ : InMux
    port map (
            O => \N__37301\,
            I => \N__37297\
        );

    \I__8076\ : InMux
    port map (
            O => \N__37300\,
            I => \N__37294\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__37297\,
            I => \N__37291\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__37294\,
            I => \N__37287\
        );

    \I__8073\ : Span4Mux_h
    port map (
            O => \N__37291\,
            I => \N__37284\
        );

    \I__8072\ : InMux
    port map (
            O => \N__37290\,
            I => \N__37281\
        );

    \I__8071\ : Odrv4
    port map (
            O => \N__37287\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__8070\ : Odrv4
    port map (
            O => \N__37284\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__37281\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__8068\ : InMux
    port map (
            O => \N__37274\,
            I => \N__37271\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__37271\,
            I => \N__37267\
        );

    \I__8066\ : InMux
    port map (
            O => \N__37270\,
            I => \N__37264\
        );

    \I__8065\ : Odrv12
    port map (
            O => \N__37267\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__37264\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8063\ : InMux
    port map (
            O => \N__37259\,
            I => \N__37255\
        );

    \I__8062\ : InMux
    port map (
            O => \N__37258\,
            I => \N__37252\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__37255\,
            I => \N__37249\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__37252\,
            I => \N__37246\
        );

    \I__8059\ : Span4Mux_v
    port map (
            O => \N__37249\,
            I => \N__37240\
        );

    \I__8058\ : Span4Mux_v
    port map (
            O => \N__37246\,
            I => \N__37240\
        );

    \I__8057\ : InMux
    port map (
            O => \N__37245\,
            I => \N__37237\
        );

    \I__8056\ : Odrv4
    port map (
            O => \N__37240\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__37237\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__8054\ : InMux
    port map (
            O => \N__37232\,
            I => \N__37229\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__37229\,
            I => \N__37225\
        );

    \I__8052\ : InMux
    port map (
            O => \N__37228\,
            I => \N__37222\
        );

    \I__8051\ : Odrv4
    port map (
            O => \N__37225\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__37222\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__8049\ : CascadeMux
    port map (
            O => \N__37217\,
            I => \N__37213\
        );

    \I__8048\ : InMux
    port map (
            O => \N__37216\,
            I => \N__37210\
        );

    \I__8047\ : InMux
    port map (
            O => \N__37213\,
            I => \N__37207\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__37210\,
            I => \N__37204\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__37207\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_1Z0Z_9\
        );

    \I__8044\ : Odrv4
    port map (
            O => \N__37204\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_1Z0Z_9\
        );

    \I__8043\ : CascadeMux
    port map (
            O => \N__37199\,
            I => \N__37196\
        );

    \I__8042\ : InMux
    port map (
            O => \N__37196\,
            I => \N__37192\
        );

    \I__8041\ : InMux
    port map (
            O => \N__37195\,
            I => \N__37189\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__37192\,
            I => \N__37186\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__37189\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9\
        );

    \I__8038\ : Odrv4
    port map (
            O => \N__37186\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9\
        );

    \I__8037\ : InMux
    port map (
            O => \N__37181\,
            I => \N__37177\
        );

    \I__8036\ : CascadeMux
    port map (
            O => \N__37180\,
            I => \N__37174\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__37177\,
            I => \N__37171\
        );

    \I__8034\ : InMux
    port map (
            O => \N__37174\,
            I => \N__37167\
        );

    \I__8033\ : Span4Mux_h
    port map (
            O => \N__37171\,
            I => \N__37164\
        );

    \I__8032\ : InMux
    port map (
            O => \N__37170\,
            I => \N__37161\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__37167\,
            I => \elapsed_time_ns_1_RNIAE2591_0_2\
        );

    \I__8030\ : Odrv4
    port map (
            O => \N__37164\,
            I => \elapsed_time_ns_1_RNIAE2591_0_2\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__37161\,
            I => \elapsed_time_ns_1_RNIAE2591_0_2\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__37154\,
            I => \N__37150\
        );

    \I__8027\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37147\
        );

    \I__8026\ : InMux
    port map (
            O => \N__37150\,
            I => \N__37143\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__37147\,
            I => \N__37140\
        );

    \I__8024\ : InMux
    port map (
            O => \N__37146\,
            I => \N__37137\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__37143\,
            I => \N__37134\
        );

    \I__8022\ : Odrv4
    port map (
            O => \N__37140\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_0_2\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__37137\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_0_2\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__37134\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_0_2\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__37127\,
            I => \N__37124\
        );

    \I__8018\ : InMux
    port map (
            O => \N__37124\,
            I => \N__37121\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__37121\,
            I => \N__37117\
        );

    \I__8016\ : CascadeMux
    port map (
            O => \N__37120\,
            I => \N__37114\
        );

    \I__8015\ : Span4Mux_v
    port map (
            O => \N__37117\,
            I => \N__37109\
        );

    \I__8014\ : InMux
    port map (
            O => \N__37114\,
            I => \N__37106\
        );

    \I__8013\ : InMux
    port map (
            O => \N__37113\,
            I => \N__37103\
        );

    \I__8012\ : InMux
    port map (
            O => \N__37112\,
            I => \N__37100\
        );

    \I__8011\ : Odrv4
    port map (
            O => \N__37109\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__37106\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__37103\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__37100\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2\
        );

    \I__8007\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37088\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__37088\,
            I => \N__37083\
        );

    \I__8005\ : InMux
    port map (
            O => \N__37087\,
            I => \N__37080\
        );

    \I__8004\ : InMux
    port map (
            O => \N__37086\,
            I => \N__37075\
        );

    \I__8003\ : Span12Mux_v
    port map (
            O => \N__37083\,
            I => \N__37070\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__37080\,
            I => \N__37070\
        );

    \I__8001\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37067\
        );

    \I__8000\ : InMux
    port map (
            O => \N__37078\,
            I => \N__37064\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__37075\,
            I => \N__37061\
        );

    \I__7998\ : Span12Mux_s11_h
    port map (
            O => \N__37070\,
            I => \N__37056\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__37067\,
            I => \N__37056\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__37064\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__7995\ : Odrv4
    port map (
            O => \N__37061\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__7994\ : Odrv12
    port map (
            O => \N__37056\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__7993\ : CascadeMux
    port map (
            O => \N__37049\,
            I => \N__37046\
        );

    \I__7992\ : InMux
    port map (
            O => \N__37046\,
            I => \N__37043\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__37043\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2\
        );

    \I__7990\ : CascadeMux
    port map (
            O => \N__37040\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2_cascade_\
        );

    \I__7989\ : CascadeMux
    port map (
            O => \N__37037\,
            I => \N__37034\
        );

    \I__7988\ : InMux
    port map (
            O => \N__37034\,
            I => \N__37030\
        );

    \I__7987\ : CascadeMux
    port map (
            O => \N__37033\,
            I => \N__37026\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__37030\,
            I => \N__37023\
        );

    \I__7985\ : CascadeMux
    port map (
            O => \N__37029\,
            I => \N__37015\
        );

    \I__7984\ : InMux
    port map (
            O => \N__37026\,
            I => \N__37012\
        );

    \I__7983\ : Span4Mux_h
    port map (
            O => \N__37023\,
            I => \N__37009\
        );

    \I__7982\ : InMux
    port map (
            O => \N__37022\,
            I => \N__37006\
        );

    \I__7981\ : InMux
    port map (
            O => \N__37021\,
            I => \N__37003\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37020\,
            I => \N__37000\
        );

    \I__7979\ : InMux
    port map (
            O => \N__37019\,
            I => \N__36995\
        );

    \I__7978\ : InMux
    port map (
            O => \N__37018\,
            I => \N__36995\
        );

    \I__7977\ : InMux
    port map (
            O => \N__37015\,
            I => \N__36992\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__37012\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7975\ : Odrv4
    port map (
            O => \N__37009\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__37006\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__37003\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__37000\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__36995\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__36992\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7969\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36974\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__36974\,
            I => \N__36971\
        );

    \I__7967\ : Span4Mux_h
    port map (
            O => \N__36971\,
            I => \N__36965\
        );

    \I__7966\ : InMux
    port map (
            O => \N__36970\,
            I => \N__36962\
        );

    \I__7965\ : InMux
    port map (
            O => \N__36969\,
            I => \N__36959\
        );

    \I__7964\ : InMux
    port map (
            O => \N__36968\,
            I => \N__36956\
        );

    \I__7963\ : Odrv4
    port map (
            O => \N__36965\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__36962\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__36959\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__36956\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9\
        );

    \I__7959\ : InMux
    port map (
            O => \N__36947\,
            I => \N__36944\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__36944\,
            I => \N__36939\
        );

    \I__7957\ : InMux
    port map (
            O => \N__36943\,
            I => \N__36936\
        );

    \I__7956\ : InMux
    port map (
            O => \N__36942\,
            I => \N__36933\
        );

    \I__7955\ : Odrv4
    port map (
            O => \N__36939\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__36936\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__36933\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__7952\ : InMux
    port map (
            O => \N__36926\,
            I => \N__36923\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__36923\,
            I => \N__36919\
        );

    \I__7950\ : InMux
    port map (
            O => \N__36922\,
            I => \N__36914\
        );

    \I__7949\ : Span4Mux_v
    port map (
            O => \N__36919\,
            I => \N__36911\
        );

    \I__7948\ : InMux
    port map (
            O => \N__36918\,
            I => \N__36906\
        );

    \I__7947\ : InMux
    port map (
            O => \N__36917\,
            I => \N__36906\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__36914\,
            I => \elapsed_time_ns_1_RNI1OL2M1_0_9\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__36911\,
            I => \elapsed_time_ns_1_RNI1OL2M1_0_9\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__36906\,
            I => \elapsed_time_ns_1_RNI1OL2M1_0_9\
        );

    \I__7943\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36895\
        );

    \I__7942\ : InMux
    port map (
            O => \N__36898\,
            I => \N__36892\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__36895\,
            I => \phase_controller_inst1.stoper_tr.N_244\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__36892\,
            I => \phase_controller_inst1.stoper_tr.N_244\
        );

    \I__7939\ : InMux
    port map (
            O => \N__36887\,
            I => \N__36884\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__36884\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_0_6\
        );

    \I__7937\ : CascadeMux
    port map (
            O => \N__36881\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9_cascade_\
        );

    \I__7936\ : CascadeMux
    port map (
            O => \N__36878\,
            I => \phase_controller_inst1.stoper_tr.N_249_cascade_\
        );

    \I__7935\ : CascadeMux
    port map (
            O => \N__36875\,
            I => \N__36872\
        );

    \I__7934\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36868\
        );

    \I__7933\ : InMux
    port map (
            O => \N__36871\,
            I => \N__36864\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36861\
        );

    \I__7931\ : CascadeMux
    port map (
            O => \N__36867\,
            I => \N__36858\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__36864\,
            I => \N__36855\
        );

    \I__7929\ : Span4Mux_h
    port map (
            O => \N__36861\,
            I => \N__36852\
        );

    \I__7928\ : InMux
    port map (
            O => \N__36858\,
            I => \N__36849\
        );

    \I__7927\ : Odrv4
    port map (
            O => \N__36855\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__7926\ : Odrv4
    port map (
            O => \N__36852\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__36849\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__7924\ : InMux
    port map (
            O => \N__36842\,
            I => \N__36838\
        );

    \I__7923\ : InMux
    port map (
            O => \N__36841\,
            I => \N__36833\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__36838\,
            I => \N__36830\
        );

    \I__7921\ : InMux
    port map (
            O => \N__36837\,
            I => \N__36827\
        );

    \I__7920\ : InMux
    port map (
            O => \N__36836\,
            I => \N__36824\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__36833\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__7918\ : Odrv4
    port map (
            O => \N__36830\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__36827\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__36824\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__7915\ : InMux
    port map (
            O => \N__36815\,
            I => \N__36810\
        );

    \I__7914\ : InMux
    port map (
            O => \N__36814\,
            I => \N__36807\
        );

    \I__7913\ : InMux
    port map (
            O => \N__36813\,
            I => \N__36804\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__36810\,
            I => \N__36801\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__36807\,
            I => \N__36798\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__36804\,
            I => \N__36795\
        );

    \I__7909\ : Span4Mux_h
    port map (
            O => \N__36801\,
            I => \N__36789\
        );

    \I__7908\ : Span4Mux_h
    port map (
            O => \N__36798\,
            I => \N__36789\
        );

    \I__7907\ : Span4Mux_h
    port map (
            O => \N__36795\,
            I => \N__36786\
        );

    \I__7906\ : InMux
    port map (
            O => \N__36794\,
            I => \N__36783\
        );

    \I__7905\ : Odrv4
    port map (
            O => \N__36789\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6\
        );

    \I__7904\ : Odrv4
    port map (
            O => \N__36786\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__36783\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6\
        );

    \I__7902\ : InMux
    port map (
            O => \N__36776\,
            I => \N__36771\
        );

    \I__7901\ : CascadeMux
    port map (
            O => \N__36775\,
            I => \N__36767\
        );

    \I__7900\ : InMux
    port map (
            O => \N__36774\,
            I => \N__36764\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__36771\,
            I => \N__36761\
        );

    \I__7898\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36758\
        );

    \I__7897\ : InMux
    port map (
            O => \N__36767\,
            I => \N__36755\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__36764\,
            I => \N__36752\
        );

    \I__7895\ : Span4Mux_h
    port map (
            O => \N__36761\,
            I => \N__36748\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__36758\,
            I => \N__36743\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__36755\,
            I => \N__36743\
        );

    \I__7892\ : Span4Mux_h
    port map (
            O => \N__36752\,
            I => \N__36740\
        );

    \I__7891\ : InMux
    port map (
            O => \N__36751\,
            I => \N__36737\
        );

    \I__7890\ : Odrv4
    port map (
            O => \N__36748\,
            I => \phase_controller_inst1.stoper_tr.N_250\
        );

    \I__7889\ : Odrv12
    port map (
            O => \N__36743\,
            I => \phase_controller_inst1.stoper_tr.N_250\
        );

    \I__7888\ : Odrv4
    port map (
            O => \N__36740\,
            I => \phase_controller_inst1.stoper_tr.N_250\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__36737\,
            I => \phase_controller_inst1.stoper_tr.N_250\
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__36728\,
            I => \N__36725\
        );

    \I__7885\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36719\
        );

    \I__7884\ : InMux
    port map (
            O => \N__36724\,
            I => \N__36719\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__36719\,
            I => \N__36716\
        );

    \I__7882\ : Span4Mux_v
    port map (
            O => \N__36716\,
            I => \N__36711\
        );

    \I__7881\ : InMux
    port map (
            O => \N__36715\,
            I => \N__36706\
        );

    \I__7880\ : InMux
    port map (
            O => \N__36714\,
            I => \N__36706\
        );

    \I__7879\ : Span4Mux_v
    port map (
            O => \N__36711\,
            I => \N__36703\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__36706\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7877\ : Odrv4
    port map (
            O => \N__36703\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7876\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36693\
        );

    \I__7875\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36687\
        );

    \I__7874\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36687\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__36693\,
            I => \N__36684\
        );

    \I__7872\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36681\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__36687\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7870\ : Odrv4
    port map (
            O => \N__36684\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__36681\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7868\ : InMux
    port map (
            O => \N__36674\,
            I => \N__36665\
        );

    \I__7867\ : InMux
    port map (
            O => \N__36673\,
            I => \N__36665\
        );

    \I__7866\ : InMux
    port map (
            O => \N__36672\,
            I => \N__36665\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__36665\,
            I => \N__36662\
        );

    \I__7864\ : Span4Mux_v
    port map (
            O => \N__36662\,
            I => \N__36659\
        );

    \I__7863\ : Span4Mux_v
    port map (
            O => \N__36659\,
            I => \N__36656\
        );

    \I__7862\ : Odrv4
    port map (
            O => \N__36656\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7861\ : IoInMux
    port map (
            O => \N__36653\,
            I => \N__36650\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__36650\,
            I => \N__36647\
        );

    \I__7859\ : Span4Mux_s0_v
    port map (
            O => \N__36647\,
            I => \N__36644\
        );

    \I__7858\ : Span4Mux_h
    port map (
            O => \N__36644\,
            I => \N__36641\
        );

    \I__7857\ : Span4Mux_v
    port map (
            O => \N__36641\,
            I => \N__36638\
        );

    \I__7856\ : Span4Mux_v
    port map (
            O => \N__36638\,
            I => \N__36635\
        );

    \I__7855\ : Odrv4
    port map (
            O => \N__36635\,
            I => \delay_measurement_inst.delay_tr_timer.N_434_i\
        );

    \I__7854\ : CascadeMux
    port map (
            O => \N__36632\,
            I => \N__36627\
        );

    \I__7853\ : InMux
    port map (
            O => \N__36631\,
            I => \N__36624\
        );

    \I__7852\ : InMux
    port map (
            O => \N__36630\,
            I => \N__36620\
        );

    \I__7851\ : InMux
    port map (
            O => \N__36627\,
            I => \N__36617\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__36624\,
            I => \N__36614\
        );

    \I__7849\ : InMux
    port map (
            O => \N__36623\,
            I => \N__36611\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__36620\,
            I => \N__36606\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__36617\,
            I => \N__36606\
        );

    \I__7846\ : Span12Mux_h
    port map (
            O => \N__36614\,
            I => \N__36603\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__36611\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__7844\ : Odrv12
    port map (
            O => \N__36606\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__7843\ : Odrv12
    port map (
            O => \N__36603\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__7842\ : InMux
    port map (
            O => \N__36596\,
            I => \N__36593\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__36593\,
            I => \N__36590\
        );

    \I__7840\ : Span4Mux_v
    port map (
            O => \N__36590\,
            I => \N__36585\
        );

    \I__7839\ : InMux
    port map (
            O => \N__36589\,
            I => \N__36580\
        );

    \I__7838\ : InMux
    port map (
            O => \N__36588\,
            I => \N__36580\
        );

    \I__7837\ : Span4Mux_h
    port map (
            O => \N__36585\,
            I => \N__36577\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__36580\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7835\ : Odrv4
    port map (
            O => \N__36577\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7834\ : InMux
    port map (
            O => \N__36572\,
            I => \N__36569\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__36569\,
            I => \N__36566\
        );

    \I__7832\ : Span4Mux_h
    port map (
            O => \N__36566\,
            I => \N__36563\
        );

    \I__7831\ : Span4Mux_h
    port map (
            O => \N__36563\,
            I => \N__36560\
        );

    \I__7830\ : Span4Mux_v
    port map (
            O => \N__36560\,
            I => \N__36557\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__36557\,
            I => \phase_controller_inst1.N_55\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__36554\,
            I => \N__36550\
        );

    \I__7827\ : InMux
    port map (
            O => \N__36553\,
            I => \N__36544\
        );

    \I__7826\ : InMux
    port map (
            O => \N__36550\,
            I => \N__36534\
        );

    \I__7825\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36534\
        );

    \I__7824\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36531\
        );

    \I__7823\ : CascadeMux
    port map (
            O => \N__36547\,
            I => \N__36526\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__36544\,
            I => \N__36521\
        );

    \I__7821\ : CascadeMux
    port map (
            O => \N__36543\,
            I => \N__36503\
        );

    \I__7820\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36493\
        );

    \I__7819\ : InMux
    port map (
            O => \N__36541\,
            I => \N__36493\
        );

    \I__7818\ : InMux
    port map (
            O => \N__36540\,
            I => \N__36493\
        );

    \I__7817\ : InMux
    port map (
            O => \N__36539\,
            I => \N__36493\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__36534\,
            I => \N__36488\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__36531\,
            I => \N__36488\
        );

    \I__7814\ : InMux
    port map (
            O => \N__36530\,
            I => \N__36485\
        );

    \I__7813\ : InMux
    port map (
            O => \N__36529\,
            I => \N__36480\
        );

    \I__7812\ : InMux
    port map (
            O => \N__36526\,
            I => \N__36480\
        );

    \I__7811\ : InMux
    port map (
            O => \N__36525\,
            I => \N__36477\
        );

    \I__7810\ : InMux
    port map (
            O => \N__36524\,
            I => \N__36474\
        );

    \I__7809\ : Span4Mux_v
    port map (
            O => \N__36521\,
            I => \N__36471\
        );

    \I__7808\ : InMux
    port map (
            O => \N__36520\,
            I => \N__36466\
        );

    \I__7807\ : InMux
    port map (
            O => \N__36519\,
            I => \N__36466\
        );

    \I__7806\ : InMux
    port map (
            O => \N__36518\,
            I => \N__36459\
        );

    \I__7805\ : InMux
    port map (
            O => \N__36517\,
            I => \N__36459\
        );

    \I__7804\ : InMux
    port map (
            O => \N__36516\,
            I => \N__36459\
        );

    \I__7803\ : InMux
    port map (
            O => \N__36515\,
            I => \N__36454\
        );

    \I__7802\ : InMux
    port map (
            O => \N__36514\,
            I => \N__36454\
        );

    \I__7801\ : InMux
    port map (
            O => \N__36513\,
            I => \N__36443\
        );

    \I__7800\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36443\
        );

    \I__7799\ : InMux
    port map (
            O => \N__36511\,
            I => \N__36443\
        );

    \I__7798\ : InMux
    port map (
            O => \N__36510\,
            I => \N__36443\
        );

    \I__7797\ : InMux
    port map (
            O => \N__36509\,
            I => \N__36443\
        );

    \I__7796\ : InMux
    port map (
            O => \N__36508\,
            I => \N__36434\
        );

    \I__7795\ : InMux
    port map (
            O => \N__36507\,
            I => \N__36434\
        );

    \I__7794\ : InMux
    port map (
            O => \N__36506\,
            I => \N__36434\
        );

    \I__7793\ : InMux
    port map (
            O => \N__36503\,
            I => \N__36434\
        );

    \I__7792\ : InMux
    port map (
            O => \N__36502\,
            I => \N__36431\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__36493\,
            I => \N__36426\
        );

    \I__7790\ : Span4Mux_h
    port map (
            O => \N__36488\,
            I => \N__36426\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__36485\,
            I => \N__36421\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__36480\,
            I => \N__36421\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__36477\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__36474\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7785\ : Odrv4
    port map (
            O => \N__36471\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__36466\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__36459\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__36454\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__36443\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__36434\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__36431\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7778\ : Odrv4
    port map (
            O => \N__36426\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7777\ : Odrv4
    port map (
            O => \N__36421\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__7776\ : CascadeMux
    port map (
            O => \N__36398\,
            I => \N__36393\
        );

    \I__7775\ : CascadeMux
    port map (
            O => \N__36397\,
            I => \N__36390\
        );

    \I__7774\ : CascadeMux
    port map (
            O => \N__36396\,
            I => \N__36386\
        );

    \I__7773\ : InMux
    port map (
            O => \N__36393\,
            I => \N__36378\
        );

    \I__7772\ : InMux
    port map (
            O => \N__36390\,
            I => \N__36378\
        );

    \I__7771\ : InMux
    port map (
            O => \N__36389\,
            I => \N__36378\
        );

    \I__7770\ : InMux
    port map (
            O => \N__36386\,
            I => \N__36371\
        );

    \I__7769\ : InMux
    port map (
            O => \N__36385\,
            I => \N__36371\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__36378\,
            I => \N__36367\
        );

    \I__7767\ : InMux
    port map (
            O => \N__36377\,
            I => \N__36364\
        );

    \I__7766\ : CascadeMux
    port map (
            O => \N__36376\,
            I => \N__36359\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__36371\,
            I => \N__36356\
        );

    \I__7764\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36353\
        );

    \I__7763\ : Span4Mux_v
    port map (
            O => \N__36367\,
            I => \N__36348\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__36364\,
            I => \N__36348\
        );

    \I__7761\ : InMux
    port map (
            O => \N__36363\,
            I => \N__36343\
        );

    \I__7760\ : InMux
    port map (
            O => \N__36362\,
            I => \N__36343\
        );

    \I__7759\ : InMux
    port map (
            O => \N__36359\,
            I => \N__36340\
        );

    \I__7758\ : Odrv4
    port map (
            O => \N__36356\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__36353\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__7756\ : Odrv4
    port map (
            O => \N__36348\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__36343\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__36340\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__7753\ : CascadeMux
    port map (
            O => \N__36329\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_\
        );

    \I__7752\ : InMux
    port map (
            O => \N__36326\,
            I => \N__36323\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__36323\,
            I => \N__36318\
        );

    \I__7750\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36315\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__36321\,
            I => \N__36311\
        );

    \I__7748\ : Span4Mux_v
    port map (
            O => \N__36318\,
            I => \N__36304\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__36315\,
            I => \N__36301\
        );

    \I__7746\ : InMux
    port map (
            O => \N__36314\,
            I => \N__36298\
        );

    \I__7745\ : InMux
    port map (
            O => \N__36311\,
            I => \N__36293\
        );

    \I__7744\ : InMux
    port map (
            O => \N__36310\,
            I => \N__36293\
        );

    \I__7743\ : InMux
    port map (
            O => \N__36309\,
            I => \N__36288\
        );

    \I__7742\ : InMux
    port map (
            O => \N__36308\,
            I => \N__36288\
        );

    \I__7741\ : InMux
    port map (
            O => \N__36307\,
            I => \N__36285\
        );

    \I__7740\ : Span4Mux_h
    port map (
            O => \N__36304\,
            I => \N__36282\
        );

    \I__7739\ : Odrv4
    port map (
            O => \N__36301\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__36298\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__36293\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__36288\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__36285\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__7734\ : Odrv4
    port map (
            O => \N__36282\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__7733\ : CascadeMux
    port map (
            O => \N__36269\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_\
        );

    \I__7732\ : InMux
    port map (
            O => \N__36266\,
            I => \N__36261\
        );

    \I__7731\ : InMux
    port map (
            O => \N__36265\,
            I => \N__36256\
        );

    \I__7730\ : InMux
    port map (
            O => \N__36264\,
            I => \N__36256\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__36261\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__36256\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\
        );

    \I__7727\ : InMux
    port map (
            O => \N__36251\,
            I => \N__36244\
        );

    \I__7726\ : InMux
    port map (
            O => \N__36250\,
            I => \N__36244\
        );

    \I__7725\ : InMux
    port map (
            O => \N__36249\,
            I => \N__36241\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__36244\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__36241\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\
        );

    \I__7722\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36233\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__36233\,
            I => \N__36229\
        );

    \I__7720\ : InMux
    port map (
            O => \N__36232\,
            I => \N__36226\
        );

    \I__7719\ : Odrv4
    port map (
            O => \N__36229\,
            I => \elapsed_time_ns_1_RNI0GIF91_0_26\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__36226\,
            I => \elapsed_time_ns_1_RNI0GIF91_0_26\
        );

    \I__7717\ : InMux
    port map (
            O => \N__36221\,
            I => \N__36218\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__36218\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6\
        );

    \I__7715\ : CascadeMux
    port map (
            O => \N__36215\,
            I => \N__36212\
        );

    \I__7714\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36209\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__36209\,
            I => \elapsed_time_ns_1_RNITCIF91_0_23\
        );

    \I__7712\ : CascadeMux
    port map (
            O => \N__36206\,
            I => \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\
        );

    \I__7711\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36200\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__36200\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_0_15\
        );

    \I__7709\ : CascadeMux
    port map (
            O => \N__36197\,
            I => \N__36194\
        );

    \I__7708\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36190\
        );

    \I__7707\ : InMux
    port map (
            O => \N__36193\,
            I => \N__36187\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__36190\,
            I => \elapsed_time_ns_1_RNI1HIF91_0_27\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__36187\,
            I => \elapsed_time_ns_1_RNI1HIF91_0_27\
        );

    \I__7704\ : InMux
    port map (
            O => \N__36182\,
            I => \N__36179\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__36179\,
            I => \N__36173\
        );

    \I__7702\ : CascadeMux
    port map (
            O => \N__36178\,
            I => \N__36168\
        );

    \I__7701\ : CascadeMux
    port map (
            O => \N__36177\,
            I => \N__36164\
        );

    \I__7700\ : CascadeMux
    port map (
            O => \N__36176\,
            I => \N__36160\
        );

    \I__7699\ : Span4Mux_h
    port map (
            O => \N__36173\,
            I => \N__36157\
        );

    \I__7698\ : CascadeMux
    port map (
            O => \N__36172\,
            I => \N__36149\
        );

    \I__7697\ : CascadeMux
    port map (
            O => \N__36171\,
            I => \N__36146\
        );

    \I__7696\ : InMux
    port map (
            O => \N__36168\,
            I => \N__36141\
        );

    \I__7695\ : InMux
    port map (
            O => \N__36167\,
            I => \N__36138\
        );

    \I__7694\ : InMux
    port map (
            O => \N__36164\,
            I => \N__36135\
        );

    \I__7693\ : InMux
    port map (
            O => \N__36163\,
            I => \N__36130\
        );

    \I__7692\ : InMux
    port map (
            O => \N__36160\,
            I => \N__36130\
        );

    \I__7691\ : Span4Mux_v
    port map (
            O => \N__36157\,
            I => \N__36121\
        );

    \I__7690\ : InMux
    port map (
            O => \N__36156\,
            I => \N__36114\
        );

    \I__7689\ : InMux
    port map (
            O => \N__36155\,
            I => \N__36114\
        );

    \I__7688\ : InMux
    port map (
            O => \N__36154\,
            I => \N__36114\
        );

    \I__7687\ : InMux
    port map (
            O => \N__36153\,
            I => \N__36107\
        );

    \I__7686\ : InMux
    port map (
            O => \N__36152\,
            I => \N__36107\
        );

    \I__7685\ : InMux
    port map (
            O => \N__36149\,
            I => \N__36107\
        );

    \I__7684\ : InMux
    port map (
            O => \N__36146\,
            I => \N__36100\
        );

    \I__7683\ : InMux
    port map (
            O => \N__36145\,
            I => \N__36100\
        );

    \I__7682\ : InMux
    port map (
            O => \N__36144\,
            I => \N__36100\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__36141\,
            I => \N__36091\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__36138\,
            I => \N__36091\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__36135\,
            I => \N__36091\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__36130\,
            I => \N__36091\
        );

    \I__7677\ : InMux
    port map (
            O => \N__36129\,
            I => \N__36088\
        );

    \I__7676\ : InMux
    port map (
            O => \N__36128\,
            I => \N__36081\
        );

    \I__7675\ : InMux
    port map (
            O => \N__36127\,
            I => \N__36081\
        );

    \I__7674\ : InMux
    port map (
            O => \N__36126\,
            I => \N__36081\
        );

    \I__7673\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36076\
        );

    \I__7672\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36076\
        );

    \I__7671\ : Odrv4
    port map (
            O => \N__36121\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__36114\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__36107\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__36100\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__7667\ : Odrv4
    port map (
            O => \N__36091\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__36088\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__36081\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__36076\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__7663\ : CascadeMux
    port map (
            O => \N__36059\,
            I => \N__36056\
        );

    \I__7662\ : InMux
    port map (
            O => \N__36056\,
            I => \N__36052\
        );

    \I__7661\ : InMux
    port map (
            O => \N__36055\,
            I => \N__36049\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__36052\,
            I => \elapsed_time_ns_1_RNIUDIF91_0_24\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__36049\,
            I => \elapsed_time_ns_1_RNIUDIF91_0_24\
        );

    \I__7658\ : CascadeMux
    port map (
            O => \N__36044\,
            I => \delay_measurement_inst.delay_tr_timer.N_367_cascade_\
        );

    \I__7657\ : InMux
    port map (
            O => \N__36041\,
            I => \N__36037\
        );

    \I__7656\ : InMux
    port map (
            O => \N__36040\,
            I => \N__36033\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__36037\,
            I => \N__36030\
        );

    \I__7654\ : InMux
    port map (
            O => \N__36036\,
            I => \N__36027\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__36033\,
            I => \N__36020\
        );

    \I__7652\ : Span4Mux_h
    port map (
            O => \N__36030\,
            I => \N__36020\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__36027\,
            I => \N__36020\
        );

    \I__7650\ : Odrv4
    port map (
            O => \N__36020\,
            I => \delay_measurement_inst.delay_tr_timer.N_378\
        );

    \I__7649\ : InMux
    port map (
            O => \N__36017\,
            I => \N__36014\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__36014\,
            I => \N__36011\
        );

    \I__7647\ : Span12Mux_v
    port map (
            O => \N__36011\,
            I => \N__36006\
        );

    \I__7646\ : InMux
    port map (
            O => \N__36010\,
            I => \N__36001\
        );

    \I__7645\ : InMux
    port map (
            O => \N__36009\,
            I => \N__36001\
        );

    \I__7644\ : Odrv12
    port map (
            O => \N__36006\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__36001\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__7642\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35993\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__35993\,
            I => \delay_measurement_inst.delay_tr_timer.N_349\
        );

    \I__7640\ : InMux
    port map (
            O => \N__35990\,
            I => \N__35987\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__35987\,
            I => \elapsed_time_ns_1_RNIVEIF91_0_25\
        );

    \I__7638\ : CascadeMux
    port map (
            O => \N__35984\,
            I => \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\
        );

    \I__7637\ : InMux
    port map (
            O => \N__35981\,
            I => \N__35978\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__35978\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_o5_6Z0Z_15\
        );

    \I__7635\ : CascadeMux
    port map (
            O => \N__35975\,
            I => \N__35972\
        );

    \I__7634\ : InMux
    port map (
            O => \N__35972\,
            I => \N__35968\
        );

    \I__7633\ : InMux
    port map (
            O => \N__35971\,
            I => \N__35965\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__35968\,
            I => \elapsed_time_ns_1_RNI2IIF91_0_28\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__35965\,
            I => \elapsed_time_ns_1_RNI2IIF91_0_28\
        );

    \I__7630\ : CascadeMux
    port map (
            O => \N__35960\,
            I => \N__35957\
        );

    \I__7629\ : InMux
    port map (
            O => \N__35957\,
            I => \N__35954\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__35954\,
            I => \N__35951\
        );

    \I__7627\ : Span4Mux_v
    port map (
            O => \N__35951\,
            I => \N__35947\
        );

    \I__7626\ : InMux
    port map (
            O => \N__35950\,
            I => \N__35944\
        );

    \I__7625\ : Odrv4
    port map (
            O => \N__35947\,
            I => \delay_measurement_inst.delay_tr_timer.N_345\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__35944\,
            I => \delay_measurement_inst.delay_tr_timer.N_345\
        );

    \I__7623\ : InMux
    port map (
            O => \N__35939\,
            I => \N__35936\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__35936\,
            I => \delay_measurement_inst.delay_tr_timer.N_348\
        );

    \I__7621\ : InMux
    port map (
            O => \N__35933\,
            I => \N__35930\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__35930\,
            I => \delay_measurement_inst.delay_tr_timer.N_347\
        );

    \I__7619\ : CascadeMux
    port map (
            O => \N__35927\,
            I => \delay_measurement_inst.delay_tr_timer.N_347_cascade_\
        );

    \I__7618\ : CascadeMux
    port map (
            O => \N__35924\,
            I => \N__35921\
        );

    \I__7617\ : InMux
    port map (
            O => \N__35921\,
            I => \N__35915\
        );

    \I__7616\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35915\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__35915\,
            I => \N__35911\
        );

    \I__7614\ : InMux
    port map (
            O => \N__35914\,
            I => \N__35908\
        );

    \I__7613\ : Span4Mux_h
    port map (
            O => \N__35911\,
            I => \N__35905\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__35908\,
            I => \delay_measurement_inst.delay_tr_timer.N_365\
        );

    \I__7611\ : Odrv4
    port map (
            O => \N__35905\,
            I => \delay_measurement_inst.delay_tr_timer.N_365\
        );

    \I__7610\ : InMux
    port map (
            O => \N__35900\,
            I => \N__35897\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__35897\,
            I => \N__35894\
        );

    \I__7608\ : Odrv4
    port map (
            O => \N__35894\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__7607\ : InMux
    port map (
            O => \N__35891\,
            I => \N__35888\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__35888\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__7605\ : CascadeMux
    port map (
            O => \N__35885\,
            I => \N__35882\
        );

    \I__7604\ : InMux
    port map (
            O => \N__35882\,
            I => \N__35879\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__35879\,
            I => \N__35874\
        );

    \I__7602\ : InMux
    port map (
            O => \N__35878\,
            I => \N__35871\
        );

    \I__7601\ : CascadeMux
    port map (
            O => \N__35877\,
            I => \N__35868\
        );

    \I__7600\ : Span4Mux_h
    port map (
            O => \N__35874\,
            I => \N__35864\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__35871\,
            I => \N__35861\
        );

    \I__7598\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35858\
        );

    \I__7597\ : InMux
    port map (
            O => \N__35867\,
            I => \N__35855\
        );

    \I__7596\ : Span4Mux_h
    port map (
            O => \N__35864\,
            I => \N__35850\
        );

    \I__7595\ : Span4Mux_v
    port map (
            O => \N__35861\,
            I => \N__35850\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__35858\,
            I => \N__35845\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__35855\,
            I => \N__35845\
        );

    \I__7592\ : Span4Mux_v
    port map (
            O => \N__35850\,
            I => \N__35842\
        );

    \I__7591\ : Span4Mux_h
    port map (
            O => \N__35845\,
            I => \N__35839\
        );

    \I__7590\ : Odrv4
    port map (
            O => \N__35842\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__7589\ : Odrv4
    port map (
            O => \N__35839\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__7588\ : InMux
    port map (
            O => \N__35834\,
            I => \N__35822\
        );

    \I__7587\ : CascadeMux
    port map (
            O => \N__35833\,
            I => \N__35815\
        );

    \I__7586\ : InMux
    port map (
            O => \N__35832\,
            I => \N__35801\
        );

    \I__7585\ : InMux
    port map (
            O => \N__35831\,
            I => \N__35801\
        );

    \I__7584\ : InMux
    port map (
            O => \N__35830\,
            I => \N__35801\
        );

    \I__7583\ : InMux
    port map (
            O => \N__35829\,
            I => \N__35801\
        );

    \I__7582\ : InMux
    port map (
            O => \N__35828\,
            I => \N__35796\
        );

    \I__7581\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35796\
        );

    \I__7580\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35791\
        );

    \I__7579\ : InMux
    port map (
            O => \N__35825\,
            I => \N__35791\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__35822\,
            I => \N__35788\
        );

    \I__7577\ : InMux
    port map (
            O => \N__35821\,
            I => \N__35779\
        );

    \I__7576\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35779\
        );

    \I__7575\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35779\
        );

    \I__7574\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35779\
        );

    \I__7573\ : InMux
    port map (
            O => \N__35815\,
            I => \N__35767\
        );

    \I__7572\ : InMux
    port map (
            O => \N__35814\,
            I => \N__35767\
        );

    \I__7571\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35767\
        );

    \I__7570\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35767\
        );

    \I__7569\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35767\
        );

    \I__7568\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35764\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__35801\,
            I => \N__35751\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__35796\,
            I => \N__35751\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__35791\,
            I => \N__35751\
        );

    \I__7564\ : Span4Mux_v
    port map (
            O => \N__35788\,
            I => \N__35748\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__35779\,
            I => \N__35745\
        );

    \I__7562\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35742\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__35767\,
            I => \N__35731\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__35764\,
            I => \N__35731\
        );

    \I__7559\ : InMux
    port map (
            O => \N__35763\,
            I => \N__35718\
        );

    \I__7558\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35718\
        );

    \I__7557\ : InMux
    port map (
            O => \N__35761\,
            I => \N__35718\
        );

    \I__7556\ : InMux
    port map (
            O => \N__35760\,
            I => \N__35718\
        );

    \I__7555\ : InMux
    port map (
            O => \N__35759\,
            I => \N__35718\
        );

    \I__7554\ : InMux
    port map (
            O => \N__35758\,
            I => \N__35718\
        );

    \I__7553\ : Span4Mux_v
    port map (
            O => \N__35751\,
            I => \N__35715\
        );

    \I__7552\ : Sp12to4
    port map (
            O => \N__35748\,
            I => \N__35712\
        );

    \I__7551\ : Span4Mux_v
    port map (
            O => \N__35745\,
            I => \N__35707\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__35742\,
            I => \N__35707\
        );

    \I__7549\ : InMux
    port map (
            O => \N__35741\,
            I => \N__35694\
        );

    \I__7548\ : InMux
    port map (
            O => \N__35740\,
            I => \N__35694\
        );

    \I__7547\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35694\
        );

    \I__7546\ : InMux
    port map (
            O => \N__35738\,
            I => \N__35694\
        );

    \I__7545\ : InMux
    port map (
            O => \N__35737\,
            I => \N__35694\
        );

    \I__7544\ : InMux
    port map (
            O => \N__35736\,
            I => \N__35694\
        );

    \I__7543\ : Span4Mux_h
    port map (
            O => \N__35731\,
            I => \N__35691\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__35718\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7541\ : Odrv4
    port map (
            O => \N__35715\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7540\ : Odrv12
    port map (
            O => \N__35712\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7539\ : Odrv4
    port map (
            O => \N__35707\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__35694\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7537\ : Odrv4
    port map (
            O => \N__35691\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7536\ : InMux
    port map (
            O => \N__35678\,
            I => \N__35666\
        );

    \I__7535\ : InMux
    port map (
            O => \N__35677\,
            I => \N__35666\
        );

    \I__7534\ : InMux
    port map (
            O => \N__35676\,
            I => \N__35661\
        );

    \I__7533\ : InMux
    port map (
            O => \N__35675\,
            I => \N__35661\
        );

    \I__7532\ : CascadeMux
    port map (
            O => \N__35674\,
            I => \N__35658\
        );

    \I__7531\ : CascadeMux
    port map (
            O => \N__35673\,
            I => \N__35655\
        );

    \I__7530\ : CascadeMux
    port map (
            O => \N__35672\,
            I => \N__35639\
        );

    \I__7529\ : CascadeMux
    port map (
            O => \N__35671\,
            I => \N__35636\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__35666\,
            I => \N__35626\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__35661\,
            I => \N__35623\
        );

    \I__7526\ : InMux
    port map (
            O => \N__35658\,
            I => \N__35610\
        );

    \I__7525\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35610\
        );

    \I__7524\ : InMux
    port map (
            O => \N__35654\,
            I => \N__35610\
        );

    \I__7523\ : InMux
    port map (
            O => \N__35653\,
            I => \N__35610\
        );

    \I__7522\ : InMux
    port map (
            O => \N__35652\,
            I => \N__35610\
        );

    \I__7521\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35610\
        );

    \I__7520\ : InMux
    port map (
            O => \N__35650\,
            I => \N__35599\
        );

    \I__7519\ : InMux
    port map (
            O => \N__35649\,
            I => \N__35599\
        );

    \I__7518\ : InMux
    port map (
            O => \N__35648\,
            I => \N__35599\
        );

    \I__7517\ : InMux
    port map (
            O => \N__35647\,
            I => \N__35599\
        );

    \I__7516\ : InMux
    port map (
            O => \N__35646\,
            I => \N__35599\
        );

    \I__7515\ : InMux
    port map (
            O => \N__35645\,
            I => \N__35590\
        );

    \I__7514\ : InMux
    port map (
            O => \N__35644\,
            I => \N__35590\
        );

    \I__7513\ : InMux
    port map (
            O => \N__35643\,
            I => \N__35590\
        );

    \I__7512\ : InMux
    port map (
            O => \N__35642\,
            I => \N__35590\
        );

    \I__7511\ : InMux
    port map (
            O => \N__35639\,
            I => \N__35575\
        );

    \I__7510\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35575\
        );

    \I__7509\ : InMux
    port map (
            O => \N__35635\,
            I => \N__35575\
        );

    \I__7508\ : InMux
    port map (
            O => \N__35634\,
            I => \N__35575\
        );

    \I__7507\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35575\
        );

    \I__7506\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35570\
        );

    \I__7505\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35570\
        );

    \I__7504\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35565\
        );

    \I__7503\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35565\
        );

    \I__7502\ : Span4Mux_v
    port map (
            O => \N__35626\,
            I => \N__35562\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__35623\,
            I => \N__35557\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__35610\,
            I => \N__35557\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__35599\,
            I => \N__35552\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__35590\,
            I => \N__35552\
        );

    \I__7497\ : InMux
    port map (
            O => \N__35589\,
            I => \N__35543\
        );

    \I__7496\ : InMux
    port map (
            O => \N__35588\,
            I => \N__35543\
        );

    \I__7495\ : InMux
    port map (
            O => \N__35587\,
            I => \N__35543\
        );

    \I__7494\ : InMux
    port map (
            O => \N__35586\,
            I => \N__35543\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__35575\,
            I => \N__35538\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__35570\,
            I => \N__35538\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__35565\,
            I => \N__35535\
        );

    \I__7490\ : Span4Mux_h
    port map (
            O => \N__35562\,
            I => \N__35528\
        );

    \I__7489\ : Span4Mux_v
    port map (
            O => \N__35557\,
            I => \N__35528\
        );

    \I__7488\ : Span4Mux_v
    port map (
            O => \N__35552\,
            I => \N__35528\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__35543\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__7486\ : Odrv4
    port map (
            O => \N__35538\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__7485\ : Odrv4
    port map (
            O => \N__35535\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__7484\ : Odrv4
    port map (
            O => \N__35528\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__7483\ : CascadeMux
    port map (
            O => \N__35519\,
            I => \N__35501\
        );

    \I__7482\ : CascadeMux
    port map (
            O => \N__35518\,
            I => \N__35498\
        );

    \I__7481\ : CascadeMux
    port map (
            O => \N__35517\,
            I => \N__35495\
        );

    \I__7480\ : CascadeMux
    port map (
            O => \N__35516\,
            I => \N__35489\
        );

    \I__7479\ : CascadeMux
    port map (
            O => \N__35515\,
            I => \N__35486\
        );

    \I__7478\ : CascadeMux
    port map (
            O => \N__35514\,
            I => \N__35483\
        );

    \I__7477\ : CascadeMux
    port map (
            O => \N__35513\,
            I => \N__35480\
        );

    \I__7476\ : CascadeMux
    port map (
            O => \N__35512\,
            I => \N__35477\
        );

    \I__7475\ : CascadeMux
    port map (
            O => \N__35511\,
            I => \N__35472\
        );

    \I__7474\ : CascadeMux
    port map (
            O => \N__35510\,
            I => \N__35469\
        );

    \I__7473\ : CascadeMux
    port map (
            O => \N__35509\,
            I => \N__35466\
        );

    \I__7472\ : CascadeMux
    port map (
            O => \N__35508\,
            I => \N__35463\
        );

    \I__7471\ : CascadeMux
    port map (
            O => \N__35507\,
            I => \N__35459\
        );

    \I__7470\ : InMux
    port map (
            O => \N__35506\,
            I => \N__35446\
        );

    \I__7469\ : InMux
    port map (
            O => \N__35505\,
            I => \N__35446\
        );

    \I__7468\ : InMux
    port map (
            O => \N__35504\,
            I => \N__35446\
        );

    \I__7467\ : InMux
    port map (
            O => \N__35501\,
            I => \N__35446\
        );

    \I__7466\ : InMux
    port map (
            O => \N__35498\,
            I => \N__35446\
        );

    \I__7465\ : InMux
    port map (
            O => \N__35495\,
            I => \N__35446\
        );

    \I__7464\ : CascadeMux
    port map (
            O => \N__35494\,
            I => \N__35440\
        );

    \I__7463\ : CascadeMux
    port map (
            O => \N__35493\,
            I => \N__35436\
        );

    \I__7462\ : CascadeMux
    port map (
            O => \N__35492\,
            I => \N__35433\
        );

    \I__7461\ : InMux
    port map (
            O => \N__35489\,
            I => \N__35426\
        );

    \I__7460\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35426\
        );

    \I__7459\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35419\
        );

    \I__7458\ : InMux
    port map (
            O => \N__35480\,
            I => \N__35419\
        );

    \I__7457\ : InMux
    port map (
            O => \N__35477\,
            I => \N__35419\
        );

    \I__7456\ : InMux
    port map (
            O => \N__35476\,
            I => \N__35410\
        );

    \I__7455\ : InMux
    port map (
            O => \N__35475\,
            I => \N__35410\
        );

    \I__7454\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35410\
        );

    \I__7453\ : InMux
    port map (
            O => \N__35469\,
            I => \N__35410\
        );

    \I__7452\ : InMux
    port map (
            O => \N__35466\,
            I => \N__35405\
        );

    \I__7451\ : InMux
    port map (
            O => \N__35463\,
            I => \N__35405\
        );

    \I__7450\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35400\
        );

    \I__7449\ : InMux
    port map (
            O => \N__35459\,
            I => \N__35400\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__35446\,
            I => \N__35397\
        );

    \I__7447\ : InMux
    port map (
            O => \N__35445\,
            I => \N__35388\
        );

    \I__7446\ : InMux
    port map (
            O => \N__35444\,
            I => \N__35388\
        );

    \I__7445\ : InMux
    port map (
            O => \N__35443\,
            I => \N__35388\
        );

    \I__7444\ : InMux
    port map (
            O => \N__35440\,
            I => \N__35388\
        );

    \I__7443\ : InMux
    port map (
            O => \N__35439\,
            I => \N__35377\
        );

    \I__7442\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35377\
        );

    \I__7441\ : InMux
    port map (
            O => \N__35433\,
            I => \N__35377\
        );

    \I__7440\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35377\
        );

    \I__7439\ : InMux
    port map (
            O => \N__35431\,
            I => \N__35377\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__35426\,
            I => \N__35372\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__35419\,
            I => \N__35372\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__35410\,
            I => \N__35365\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__35405\,
            I => \N__35365\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__35400\,
            I => \N__35365\
        );

    \I__7433\ : Span4Mux_v
    port map (
            O => \N__35397\,
            I => \N__35360\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__35388\,
            I => \N__35360\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__35377\,
            I => \N__35355\
        );

    \I__7430\ : Span4Mux_h
    port map (
            O => \N__35372\,
            I => \N__35355\
        );

    \I__7429\ : Span4Mux_h
    port map (
            O => \N__35365\,
            I => \N__35352\
        );

    \I__7428\ : Span4Mux_h
    port map (
            O => \N__35360\,
            I => \N__35349\
        );

    \I__7427\ : Span4Mux_h
    port map (
            O => \N__35355\,
            I => \N__35346\
        );

    \I__7426\ : Odrv4
    port map (
            O => \N__35352\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__7425\ : Odrv4
    port map (
            O => \N__35349\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__35346\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__7423\ : InMux
    port map (
            O => \N__35339\,
            I => \N__35336\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__35336\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__7421\ : CascadeMux
    port map (
            O => \N__35333\,
            I => \N__35330\
        );

    \I__7420\ : InMux
    port map (
            O => \N__35330\,
            I => \N__35325\
        );

    \I__7419\ : InMux
    port map (
            O => \N__35329\,
            I => \N__35322\
        );

    \I__7418\ : CascadeMux
    port map (
            O => \N__35328\,
            I => \N__35318\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__35325\,
            I => \N__35315\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__35322\,
            I => \N__35312\
        );

    \I__7415\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35307\
        );

    \I__7414\ : InMux
    port map (
            O => \N__35318\,
            I => \N__35307\
        );

    \I__7413\ : Span4Mux_v
    port map (
            O => \N__35315\,
            I => \N__35303\
        );

    \I__7412\ : Span4Mux_v
    port map (
            O => \N__35312\,
            I => \N__35300\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__35307\,
            I => \N__35297\
        );

    \I__7410\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35294\
        );

    \I__7409\ : Span4Mux_h
    port map (
            O => \N__35303\,
            I => \N__35291\
        );

    \I__7408\ : Sp12to4
    port map (
            O => \N__35300\,
            I => \N__35286\
        );

    \I__7407\ : Span12Mux_s8_v
    port map (
            O => \N__35297\,
            I => \N__35286\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__35294\,
            I => \N__35283\
        );

    \I__7405\ : Odrv4
    port map (
            O => \N__35291\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__7404\ : Odrv12
    port map (
            O => \N__35286\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__7403\ : Odrv4
    port map (
            O => \N__35283\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__7402\ : CascadeMux
    port map (
            O => \N__35276\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\
        );

    \I__7401\ : InMux
    port map (
            O => \N__35273\,
            I => \N__35269\
        );

    \I__7400\ : InMux
    port map (
            O => \N__35272\,
            I => \N__35266\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__35269\,
            I => \N__35261\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__35266\,
            I => \N__35261\
        );

    \I__7397\ : Odrv4
    port map (
            O => \N__35261\,
            I => \delay_measurement_inst.delay_tr_timer.N_380\
        );

    \I__7396\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35255\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__35255\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\
        );

    \I__7394\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35246\
        );

    \I__7393\ : InMux
    port map (
            O => \N__35251\,
            I => \N__35246\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__35246\,
            I => \delay_measurement_inst.delay_tr_timer.N_341\
        );

    \I__7391\ : InMux
    port map (
            O => \N__35243\,
            I => \N__35240\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__35240\,
            I => \delay_measurement_inst.delay_tr_timer.N_367\
        );

    \I__7389\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35234\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__35234\,
            I => \N__35231\
        );

    \I__7387\ : Odrv4
    port map (
            O => \N__35231\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__7386\ : CascadeMux
    port map (
            O => \N__35228\,
            I => \N__35225\
        );

    \I__7385\ : InMux
    port map (
            O => \N__35225\,
            I => \N__35222\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__35222\,
            I => \N__35218\
        );

    \I__7383\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35214\
        );

    \I__7382\ : Span4Mux_v
    port map (
            O => \N__35218\,
            I => \N__35211\
        );

    \I__7381\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35208\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__35214\,
            I => \N__35203\
        );

    \I__7379\ : Span4Mux_h
    port map (
            O => \N__35211\,
            I => \N__35198\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__35208\,
            I => \N__35198\
        );

    \I__7377\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35193\
        );

    \I__7376\ : InMux
    port map (
            O => \N__35206\,
            I => \N__35193\
        );

    \I__7375\ : Span4Mux_v
    port map (
            O => \N__35203\,
            I => \N__35188\
        );

    \I__7374\ : Span4Mux_h
    port map (
            O => \N__35198\,
            I => \N__35188\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__35193\,
            I => \N__35185\
        );

    \I__7372\ : Odrv4
    port map (
            O => \N__35188\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__7371\ : Odrv4
    port map (
            O => \N__35185\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__7370\ : InMux
    port map (
            O => \N__35180\,
            I => \N__35177\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__35177\,
            I => \N__35174\
        );

    \I__7368\ : Odrv4
    port map (
            O => \N__35174\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__7367\ : CascadeMux
    port map (
            O => \N__35171\,
            I => \N__35167\
        );

    \I__7366\ : InMux
    port map (
            O => \N__35170\,
            I => \N__35163\
        );

    \I__7365\ : InMux
    port map (
            O => \N__35167\,
            I => \N__35160\
        );

    \I__7364\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35157\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__35163\,
            I => \N__35153\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__35160\,
            I => \N__35150\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__35157\,
            I => \N__35146\
        );

    \I__7360\ : InMux
    port map (
            O => \N__35156\,
            I => \N__35143\
        );

    \I__7359\ : Span4Mux_v
    port map (
            O => \N__35153\,
            I => \N__35140\
        );

    \I__7358\ : Span12Mux_h
    port map (
            O => \N__35150\,
            I => \N__35137\
        );

    \I__7357\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35134\
        );

    \I__7356\ : Span4Mux_h
    port map (
            O => \N__35146\,
            I => \N__35129\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__35143\,
            I => \N__35129\
        );

    \I__7354\ : Odrv4
    port map (
            O => \N__35140\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__7353\ : Odrv12
    port map (
            O => \N__35137\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__35134\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__7351\ : Odrv4
    port map (
            O => \N__35129\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__7350\ : InMux
    port map (
            O => \N__35120\,
            I => \N__35117\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__35117\,
            I => \N__35114\
        );

    \I__7348\ : Odrv4
    port map (
            O => \N__35114\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__7347\ : InMux
    port map (
            O => \N__35111\,
            I => \N__35107\
        );

    \I__7346\ : InMux
    port map (
            O => \N__35110\,
            I => \N__35104\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__35107\,
            I => \N__35101\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__35104\,
            I => \N__35096\
        );

    \I__7343\ : Span4Mux_h
    port map (
            O => \N__35101\,
            I => \N__35093\
        );

    \I__7342\ : InMux
    port map (
            O => \N__35100\,
            I => \N__35090\
        );

    \I__7341\ : InMux
    port map (
            O => \N__35099\,
            I => \N__35087\
        );

    \I__7340\ : Span4Mux_v
    port map (
            O => \N__35096\,
            I => \N__35080\
        );

    \I__7339\ : Span4Mux_v
    port map (
            O => \N__35093\,
            I => \N__35080\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__35090\,
            I => \N__35080\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__35087\,
            I => \N__35076\
        );

    \I__7336\ : Span4Mux_h
    port map (
            O => \N__35080\,
            I => \N__35073\
        );

    \I__7335\ : InMux
    port map (
            O => \N__35079\,
            I => \N__35070\
        );

    \I__7334\ : Odrv12
    port map (
            O => \N__35076\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__7333\ : Odrv4
    port map (
            O => \N__35073\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__35070\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__7331\ : InMux
    port map (
            O => \N__35063\,
            I => \N__35060\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__35060\,
            I => \N__35057\
        );

    \I__7329\ : Odrv4
    port map (
            O => \N__35057\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__7328\ : CascadeMux
    port map (
            O => \N__35054\,
            I => \N__35051\
        );

    \I__7327\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35048\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__35048\,
            I => \N__35044\
        );

    \I__7325\ : InMux
    port map (
            O => \N__35047\,
            I => \N__35039\
        );

    \I__7324\ : Span4Mux_v
    port map (
            O => \N__35044\,
            I => \N__35035\
        );

    \I__7323\ : InMux
    port map (
            O => \N__35043\,
            I => \N__35032\
        );

    \I__7322\ : CascadeMux
    port map (
            O => \N__35042\,
            I => \N__35029\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__35039\,
            I => \N__35026\
        );

    \I__7320\ : InMux
    port map (
            O => \N__35038\,
            I => \N__35023\
        );

    \I__7319\ : Span4Mux_h
    port map (
            O => \N__35035\,
            I => \N__35018\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__35032\,
            I => \N__35018\
        );

    \I__7317\ : InMux
    port map (
            O => \N__35029\,
            I => \N__35015\
        );

    \I__7316\ : Span4Mux_v
    port map (
            O => \N__35026\,
            I => \N__35012\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__35023\,
            I => \N__35009\
        );

    \I__7314\ : Span4Mux_h
    port map (
            O => \N__35018\,
            I => \N__35006\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__35015\,
            I => \N__35003\
        );

    \I__7312\ : Odrv4
    port map (
            O => \N__35012\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__7311\ : Odrv12
    port map (
            O => \N__35009\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__7310\ : Odrv4
    port map (
            O => \N__35006\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__7309\ : Odrv12
    port map (
            O => \N__35003\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__7308\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34990\
        );

    \I__7307\ : InMux
    port map (
            O => \N__34993\,
            I => \N__34987\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__34990\,
            I => \N__34983\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__34987\,
            I => \N__34980\
        );

    \I__7304\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34977\
        );

    \I__7303\ : Span4Mux_h
    port map (
            O => \N__34983\,
            I => \N__34974\
        );

    \I__7302\ : Span4Mux_v
    port map (
            O => \N__34980\,
            I => \N__34971\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__34977\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__7300\ : Odrv4
    port map (
            O => \N__34974\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__7299\ : Odrv4
    port map (
            O => \N__34971\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__7298\ : CascadeMux
    port map (
            O => \N__34964\,
            I => \N__34956\
        );

    \I__7297\ : CascadeMux
    port map (
            O => \N__34963\,
            I => \N__34950\
        );

    \I__7296\ : CascadeMux
    port map (
            O => \N__34962\,
            I => \N__34944\
        );

    \I__7295\ : CascadeMux
    port map (
            O => \N__34961\,
            I => \N__34939\
        );

    \I__7294\ : CascadeMux
    port map (
            O => \N__34960\,
            I => \N__34934\
        );

    \I__7293\ : CascadeMux
    port map (
            O => \N__34959\,
            I => \N__34930\
        );

    \I__7292\ : InMux
    port map (
            O => \N__34956\,
            I => \N__34927\
        );

    \I__7291\ : CascadeMux
    port map (
            O => \N__34955\,
            I => \N__34923\
        );

    \I__7290\ : CascadeMux
    port map (
            O => \N__34954\,
            I => \N__34920\
        );

    \I__7289\ : CascadeMux
    port map (
            O => \N__34953\,
            I => \N__34917\
        );

    \I__7288\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34909\
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__34949\,
            I => \N__34906\
        );

    \I__7286\ : CascadeMux
    port map (
            O => \N__34948\,
            I => \N__34902\
        );

    \I__7285\ : InMux
    port map (
            O => \N__34947\,
            I => \N__34894\
        );

    \I__7284\ : InMux
    port map (
            O => \N__34944\,
            I => \N__34891\
        );

    \I__7283\ : CascadeMux
    port map (
            O => \N__34943\,
            I => \N__34887\
        );

    \I__7282\ : InMux
    port map (
            O => \N__34942\,
            I => \N__34869\
        );

    \I__7281\ : InMux
    port map (
            O => \N__34939\,
            I => \N__34851\
        );

    \I__7280\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34851\
        );

    \I__7279\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34851\
        );

    \I__7278\ : InMux
    port map (
            O => \N__34934\,
            I => \N__34851\
        );

    \I__7277\ : InMux
    port map (
            O => \N__34933\,
            I => \N__34851\
        );

    \I__7276\ : InMux
    port map (
            O => \N__34930\,
            I => \N__34851\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__34927\,
            I => \N__34848\
        );

    \I__7274\ : InMux
    port map (
            O => \N__34926\,
            I => \N__34839\
        );

    \I__7273\ : InMux
    port map (
            O => \N__34923\,
            I => \N__34839\
        );

    \I__7272\ : InMux
    port map (
            O => \N__34920\,
            I => \N__34839\
        );

    \I__7271\ : InMux
    port map (
            O => \N__34917\,
            I => \N__34839\
        );

    \I__7270\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34834\
        );

    \I__7269\ : InMux
    port map (
            O => \N__34915\,
            I => \N__34834\
        );

    \I__7268\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34826\
        );

    \I__7267\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34826\
        );

    \I__7266\ : InMux
    port map (
            O => \N__34912\,
            I => \N__34826\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__34909\,
            I => \N__34823\
        );

    \I__7264\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34806\
        );

    \I__7263\ : InMux
    port map (
            O => \N__34905\,
            I => \N__34806\
        );

    \I__7262\ : InMux
    port map (
            O => \N__34902\,
            I => \N__34806\
        );

    \I__7261\ : InMux
    port map (
            O => \N__34901\,
            I => \N__34806\
        );

    \I__7260\ : InMux
    port map (
            O => \N__34900\,
            I => \N__34806\
        );

    \I__7259\ : InMux
    port map (
            O => \N__34899\,
            I => \N__34806\
        );

    \I__7258\ : InMux
    port map (
            O => \N__34898\,
            I => \N__34806\
        );

    \I__7257\ : InMux
    port map (
            O => \N__34897\,
            I => \N__34806\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__34894\,
            I => \N__34801\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__34891\,
            I => \N__34801\
        );

    \I__7254\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34798\
        );

    \I__7253\ : InMux
    port map (
            O => \N__34887\,
            I => \N__34787\
        );

    \I__7252\ : InMux
    port map (
            O => \N__34886\,
            I => \N__34787\
        );

    \I__7251\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34787\
        );

    \I__7250\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34787\
        );

    \I__7249\ : InMux
    port map (
            O => \N__34883\,
            I => \N__34787\
        );

    \I__7248\ : InMux
    port map (
            O => \N__34882\,
            I => \N__34782\
        );

    \I__7247\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34782\
        );

    \I__7246\ : InMux
    port map (
            O => \N__34880\,
            I => \N__34771\
        );

    \I__7245\ : InMux
    port map (
            O => \N__34879\,
            I => \N__34771\
        );

    \I__7244\ : InMux
    port map (
            O => \N__34878\,
            I => \N__34771\
        );

    \I__7243\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34771\
        );

    \I__7242\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34771\
        );

    \I__7241\ : InMux
    port map (
            O => \N__34875\,
            I => \N__34766\
        );

    \I__7240\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34766\
        );

    \I__7239\ : InMux
    port map (
            O => \N__34873\,
            I => \N__34763\
        );

    \I__7238\ : InMux
    port map (
            O => \N__34872\,
            I => \N__34760\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__34869\,
            I => \N__34757\
        );

    \I__7236\ : InMux
    port map (
            O => \N__34868\,
            I => \N__34746\
        );

    \I__7235\ : InMux
    port map (
            O => \N__34867\,
            I => \N__34746\
        );

    \I__7234\ : InMux
    port map (
            O => \N__34866\,
            I => \N__34746\
        );

    \I__7233\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34746\
        );

    \I__7232\ : InMux
    port map (
            O => \N__34864\,
            I => \N__34746\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__34851\,
            I => \N__34739\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__34848\,
            I => \N__34739\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__34839\,
            I => \N__34739\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__34834\,
            I => \N__34736\
        );

    \I__7227\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34733\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__34826\,
            I => \N__34726\
        );

    \I__7225\ : Span4Mux_v
    port map (
            O => \N__34823\,
            I => \N__34726\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__34806\,
            I => \N__34726\
        );

    \I__7223\ : Span4Mux_h
    port map (
            O => \N__34801\,
            I => \N__34711\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__34798\,
            I => \N__34711\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__34787\,
            I => \N__34711\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__34782\,
            I => \N__34711\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__34771\,
            I => \N__34711\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__34766\,
            I => \N__34711\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__34763\,
            I => \N__34711\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__34760\,
            I => \N__34708\
        );

    \I__7215\ : Span4Mux_h
    port map (
            O => \N__34757\,
            I => \N__34703\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__34746\,
            I => \N__34703\
        );

    \I__7213\ : Span4Mux_v
    port map (
            O => \N__34739\,
            I => \N__34698\
        );

    \I__7212\ : Span4Mux_v
    port map (
            O => \N__34736\,
            I => \N__34698\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__34733\,
            I => \N__34691\
        );

    \I__7210\ : Span4Mux_h
    port map (
            O => \N__34726\,
            I => \N__34691\
        );

    \I__7209\ : Span4Mux_v
    port map (
            O => \N__34711\,
            I => \N__34691\
        );

    \I__7208\ : Odrv4
    port map (
            O => \N__34708\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__34703\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7206\ : Odrv4
    port map (
            O => \N__34698\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7205\ : Odrv4
    port map (
            O => \N__34691\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7204\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34679\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__34679\,
            I => \N__34676\
        );

    \I__7202\ : Span4Mux_h
    port map (
            O => \N__34676\,
            I => \N__34673\
        );

    \I__7201\ : Odrv4
    port map (
            O => \N__34673\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_10\
        );

    \I__7200\ : CascadeMux
    port map (
            O => \N__34670\,
            I => \N__34667\
        );

    \I__7199\ : InMux
    port map (
            O => \N__34667\,
            I => \N__34664\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__34664\,
            I => \N__34661\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__34661\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\
        );

    \I__7196\ : InMux
    port map (
            O => \N__34658\,
            I => \N__34655\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__34655\,
            I => \N__34652\
        );

    \I__7194\ : Odrv4
    port map (
            O => \N__34652\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__7193\ : CascadeMux
    port map (
            O => \N__34649\,
            I => \N__34646\
        );

    \I__7192\ : InMux
    port map (
            O => \N__34646\,
            I => \N__34641\
        );

    \I__7191\ : InMux
    port map (
            O => \N__34645\,
            I => \N__34638\
        );

    \I__7190\ : InMux
    port map (
            O => \N__34644\,
            I => \N__34635\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__34641\,
            I => \N__34632\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__34638\,
            I => \N__34627\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__34635\,
            I => \N__34622\
        );

    \I__7186\ : Span4Mux_v
    port map (
            O => \N__34632\,
            I => \N__34622\
        );

    \I__7185\ : InMux
    port map (
            O => \N__34631\,
            I => \N__34619\
        );

    \I__7184\ : InMux
    port map (
            O => \N__34630\,
            I => \N__34616\
        );

    \I__7183\ : Span4Mux_v
    port map (
            O => \N__34627\,
            I => \N__34611\
        );

    \I__7182\ : Span4Mux_h
    port map (
            O => \N__34622\,
            I => \N__34611\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__34619\,
            I => \N__34608\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__34616\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__7179\ : Odrv4
    port map (
            O => \N__34611\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__34608\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__7177\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34598\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__34598\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__7175\ : CascadeMux
    port map (
            O => \N__34595\,
            I => \N__34592\
        );

    \I__7174\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34589\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__34589\,
            I => \N__34585\
        );

    \I__7172\ : CascadeMux
    port map (
            O => \N__34588\,
            I => \N__34581\
        );

    \I__7171\ : Span4Mux_v
    port map (
            O => \N__34585\,
            I => \N__34578\
        );

    \I__7170\ : InMux
    port map (
            O => \N__34584\,
            I => \N__34575\
        );

    \I__7169\ : InMux
    port map (
            O => \N__34581\,
            I => \N__34572\
        );

    \I__7168\ : Span4Mux_h
    port map (
            O => \N__34578\,
            I => \N__34567\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__34575\,
            I => \N__34567\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__34572\,
            I => \N__34563\
        );

    \I__7165\ : Span4Mux_h
    port map (
            O => \N__34567\,
            I => \N__34560\
        );

    \I__7164\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34557\
        );

    \I__7163\ : Span4Mux_h
    port map (
            O => \N__34563\,
            I => \N__34552\
        );

    \I__7162\ : Span4Mux_v
    port map (
            O => \N__34560\,
            I => \N__34552\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__34557\,
            I => \N__34549\
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__34552\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__7159\ : Odrv4
    port map (
            O => \N__34549\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__7158\ : CascadeMux
    port map (
            O => \N__34544\,
            I => \N__34541\
        );

    \I__7157\ : InMux
    port map (
            O => \N__34541\,
            I => \N__34538\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__34538\,
            I => \N__34535\
        );

    \I__7155\ : Odrv4
    port map (
            O => \N__34535\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__7154\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34529\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__34529\,
            I => \N__34524\
        );

    \I__7152\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34521\
        );

    \I__7151\ : CascadeMux
    port map (
            O => \N__34527\,
            I => \N__34518\
        );

    \I__7150\ : Span4Mux_h
    port map (
            O => \N__34524\,
            I => \N__34512\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__34521\,
            I => \N__34512\
        );

    \I__7148\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34507\
        );

    \I__7147\ : InMux
    port map (
            O => \N__34517\,
            I => \N__34507\
        );

    \I__7146\ : Span4Mux_v
    port map (
            O => \N__34512\,
            I => \N__34504\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__34507\,
            I => \N__34501\
        );

    \I__7144\ : Span4Mux_h
    port map (
            O => \N__34504\,
            I => \N__34498\
        );

    \I__7143\ : Span4Mux_h
    port map (
            O => \N__34501\,
            I => \N__34495\
        );

    \I__7142\ : Odrv4
    port map (
            O => \N__34498\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__7141\ : Odrv4
    port map (
            O => \N__34495\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__7140\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34487\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__34487\,
            I => \N__34482\
        );

    \I__7138\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34479\
        );

    \I__7137\ : InMux
    port map (
            O => \N__34485\,
            I => \N__34475\
        );

    \I__7136\ : Span4Mux_h
    port map (
            O => \N__34482\,
            I => \N__34470\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__34479\,
            I => \N__34470\
        );

    \I__7134\ : InMux
    port map (
            O => \N__34478\,
            I => \N__34467\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__34475\,
            I => \N__34464\
        );

    \I__7132\ : Span4Mux_h
    port map (
            O => \N__34470\,
            I => \N__34461\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__34467\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__7130\ : Odrv4
    port map (
            O => \N__34464\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__7129\ : Odrv4
    port map (
            O => \N__34461\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__7128\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34450\
        );

    \I__7127\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34447\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__34450\,
            I => \N__34444\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__34447\,
            I => \N__34441\
        );

    \I__7124\ : Span4Mux_h
    port map (
            O => \N__34444\,
            I => \N__34438\
        );

    \I__7123\ : Span4Mux_v
    port map (
            O => \N__34441\,
            I => \N__34432\
        );

    \I__7122\ : Span4Mux_v
    port map (
            O => \N__34438\,
            I => \N__34432\
        );

    \I__7121\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34429\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__34432\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__34429\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__7118\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34421\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__34421\,
            I => \N__34418\
        );

    \I__7116\ : Span4Mux_h
    port map (
            O => \N__34418\,
            I => \N__34415\
        );

    \I__7115\ : Span4Mux_v
    port map (
            O => \N__34415\,
            I => \N__34412\
        );

    \I__7114\ : Odrv4
    port map (
            O => \N__34412\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_6\
        );

    \I__7113\ : CascadeMux
    port map (
            O => \N__34409\,
            I => \N__34406\
        );

    \I__7112\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34403\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__34403\,
            I => \N__34400\
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__34400\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\
        );

    \I__7109\ : CascadeMux
    port map (
            O => \N__34397\,
            I => \N__34394\
        );

    \I__7108\ : InMux
    port map (
            O => \N__34394\,
            I => \N__34391\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__34391\,
            I => \N__34387\
        );

    \I__7106\ : InMux
    port map (
            O => \N__34390\,
            I => \N__34382\
        );

    \I__7105\ : Span4Mux_v
    port map (
            O => \N__34387\,
            I => \N__34378\
        );

    \I__7104\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34375\
        );

    \I__7103\ : InMux
    port map (
            O => \N__34385\,
            I => \N__34372\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__34382\,
            I => \N__34369\
        );

    \I__7101\ : InMux
    port map (
            O => \N__34381\,
            I => \N__34366\
        );

    \I__7100\ : Span4Mux_h
    port map (
            O => \N__34378\,
            I => \N__34359\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__34375\,
            I => \N__34359\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__34372\,
            I => \N__34359\
        );

    \I__7097\ : Odrv4
    port map (
            O => \N__34369\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__34366\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__7095\ : Odrv4
    port map (
            O => \N__34359\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__7094\ : InMux
    port map (
            O => \N__34352\,
            I => \N__34349\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__34349\,
            I => \current_shift_inst.PI_CTRL.integrator_i_14\
        );

    \I__7092\ : CascadeMux
    port map (
            O => \N__34346\,
            I => \N__34343\
        );

    \I__7091\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34337\
        );

    \I__7090\ : InMux
    port map (
            O => \N__34342\,
            I => \N__34334\
        );

    \I__7089\ : InMux
    port map (
            O => \N__34341\,
            I => \N__34331\
        );

    \I__7088\ : InMux
    port map (
            O => \N__34340\,
            I => \N__34328\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__34337\,
            I => \N__34325\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__34334\,
            I => \N__34321\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__34331\,
            I => \N__34316\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__34328\,
            I => \N__34316\
        );

    \I__7083\ : Span12Mux_v
    port map (
            O => \N__34325\,
            I => \N__34313\
        );

    \I__7082\ : InMux
    port map (
            O => \N__34324\,
            I => \N__34310\
        );

    \I__7081\ : Span4Mux_v
    port map (
            O => \N__34321\,
            I => \N__34307\
        );

    \I__7080\ : Span4Mux_v
    port map (
            O => \N__34316\,
            I => \N__34304\
        );

    \I__7079\ : Odrv12
    port map (
            O => \N__34313\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__34310\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7077\ : Odrv4
    port map (
            O => \N__34307\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7076\ : Odrv4
    port map (
            O => \N__34304\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7075\ : CascadeMux
    port map (
            O => \N__34295\,
            I => \N__34292\
        );

    \I__7074\ : InMux
    port map (
            O => \N__34292\,
            I => \N__34289\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__34289\,
            I => \N__34286\
        );

    \I__7072\ : Odrv4
    port map (
            O => \N__34286\,
            I => \current_shift_inst.PI_CTRL.integrator_i_19\
        );

    \I__7071\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34280\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__34280\,
            I => \N__34277\
        );

    \I__7069\ : Odrv12
    port map (
            O => \N__34277\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7\
        );

    \I__7068\ : InMux
    port map (
            O => \N__34274\,
            I => \N__34271\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__34271\,
            I => \N__34268\
        );

    \I__7066\ : Odrv4
    port map (
            O => \N__34268\,
            I => \current_shift_inst.PI_CTRL.integrator_i_24\
        );

    \I__7065\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34262\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__34262\,
            I => \current_shift_inst.PI_CTRL.integrator_i_6\
        );

    \I__7063\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34256\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__34256\,
            I => \current_shift_inst.PI_CTRL.integrator_i_10\
        );

    \I__7061\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34250\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__34250\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__7059\ : InMux
    port map (
            O => \N__34247\,
            I => \N__34244\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__34244\,
            I => \N__34241\
        );

    \I__7057\ : Span4Mux_h
    port map (
            O => \N__34241\,
            I => \N__34238\
        );

    \I__7056\ : Span4Mux_h
    port map (
            O => \N__34238\,
            I => \N__34235\
        );

    \I__7055\ : Odrv4
    port map (
            O => \N__34235\,
            I => \current_shift_inst.PI_CTRL.N_74_16\
        );

    \I__7054\ : CascadeMux
    port map (
            O => \N__34232\,
            I => \N__34229\
        );

    \I__7053\ : InMux
    port map (
            O => \N__34229\,
            I => \N__34224\
        );

    \I__7052\ : InMux
    port map (
            O => \N__34228\,
            I => \N__34219\
        );

    \I__7051\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34216\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__34224\,
            I => \N__34213\
        );

    \I__7049\ : InMux
    port map (
            O => \N__34223\,
            I => \N__34210\
        );

    \I__7048\ : InMux
    port map (
            O => \N__34222\,
            I => \N__34207\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__34219\,
            I => \N__34202\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__34216\,
            I => \N__34202\
        );

    \I__7045\ : Span4Mux_v
    port map (
            O => \N__34213\,
            I => \N__34197\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__34210\,
            I => \N__34197\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__34207\,
            I => \N__34194\
        );

    \I__7042\ : Span4Mux_v
    port map (
            O => \N__34202\,
            I => \N__34188\
        );

    \I__7041\ : Span4Mux_h
    port map (
            O => \N__34197\,
            I => \N__34188\
        );

    \I__7040\ : Span4Mux_v
    port map (
            O => \N__34194\,
            I => \N__34185\
        );

    \I__7039\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34182\
        );

    \I__7038\ : Span4Mux_h
    port map (
            O => \N__34188\,
            I => \N__34179\
        );

    \I__7037\ : Odrv4
    port map (
            O => \N__34185\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__34182\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__7035\ : Odrv4
    port map (
            O => \N__34179\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__7034\ : CascadeMux
    port map (
            O => \N__34172\,
            I => \N__34169\
        );

    \I__7033\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34166\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__34166\,
            I => \N__34163\
        );

    \I__7031\ : Odrv12
    port map (
            O => \N__34163\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\
        );

    \I__7030\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34157\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__34157\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__7028\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34151\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__34151\,
            I => \N__34148\
        );

    \I__7026\ : Odrv12
    port map (
            O => \N__34148\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__7025\ : InMux
    port map (
            O => \N__34145\,
            I => \N__34142\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__34142\,
            I => \N__34139\
        );

    \I__7023\ : Odrv12
    port map (
            O => \N__34139\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__7022\ : InMux
    port map (
            O => \N__34136\,
            I => \N__34133\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__34133\,
            I => \N__34130\
        );

    \I__7020\ : Odrv12
    port map (
            O => \N__34130\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__7019\ : InMux
    port map (
            O => \N__34127\,
            I => \N__34124\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__34124\,
            I => \N__34121\
        );

    \I__7017\ : Odrv4
    port map (
            O => \N__34121\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__7016\ : InMux
    port map (
            O => \N__34118\,
            I => \N__34115\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__34115\,
            I => \N__34112\
        );

    \I__7014\ : Odrv12
    port map (
            O => \N__34112\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__7013\ : InMux
    port map (
            O => \N__34109\,
            I => \N__34106\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__34106\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__7011\ : ClkMux
    port map (
            O => \N__34103\,
            I => \N__34100\
        );

    \I__7010\ : GlobalMux
    port map (
            O => \N__34100\,
            I => \N__34097\
        );

    \I__7009\ : gio2CtrlBuf
    port map (
            O => \N__34097\,
            I => delay_tr_input_c_g
        );

    \I__7008\ : InMux
    port map (
            O => \N__34094\,
            I => \N__34091\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__34091\,
            I => \N__34088\
        );

    \I__7006\ : Odrv4
    port map (
            O => \N__34088\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__7005\ : InMux
    port map (
            O => \N__34085\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__7004\ : InMux
    port map (
            O => \N__34082\,
            I => \N__34079\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__34079\,
            I => \N__34076\
        );

    \I__7002\ : Odrv4
    port map (
            O => \N__34076\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__7001\ : InMux
    port map (
            O => \N__34073\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__7000\ : InMux
    port map (
            O => \N__34070\,
            I => \bfn_15_20_0_\
        );

    \I__6999\ : InMux
    port map (
            O => \N__34067\,
            I => \N__34064\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__34064\,
            I => \N__34061\
        );

    \I__6997\ : Odrv4
    port map (
            O => \N__34061\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__6996\ : InMux
    port map (
            O => \N__34058\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__6995\ : InMux
    port map (
            O => \N__34055\,
            I => \N__34052\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__34052\,
            I => \N__34049\
        );

    \I__6993\ : Odrv4
    port map (
            O => \N__34049\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__6992\ : InMux
    port map (
            O => \N__34046\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__6991\ : InMux
    port map (
            O => \N__34043\,
            I => \N__34040\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__34040\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__6989\ : CascadeMux
    port map (
            O => \N__34037\,
            I => \N__34034\
        );

    \I__6988\ : InMux
    port map (
            O => \N__34034\,
            I => \N__34028\
        );

    \I__6987\ : InMux
    port map (
            O => \N__34033\,
            I => \N__34028\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__34028\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__6985\ : InMux
    port map (
            O => \N__34025\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__6984\ : InMux
    port map (
            O => \N__34022\,
            I => \N__34019\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__34019\,
            I => \N__34016\
        );

    \I__6982\ : Odrv4
    port map (
            O => \N__34016\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__6981\ : InMux
    port map (
            O => \N__34013\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__6980\ : InMux
    port map (
            O => \N__34010\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__6979\ : InMux
    port map (
            O => \N__34007\,
            I => \N__34004\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__34004\,
            I => \N__34001\
        );

    \I__6977\ : Span4Mux_h
    port map (
            O => \N__34001\,
            I => \N__33998\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__33998\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__33995\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\
        );

    \I__6974\ : InMux
    port map (
            O => \N__33992\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__6973\ : InMux
    port map (
            O => \N__33989\,
            I => \N__33986\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__33986\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__6971\ : InMux
    port map (
            O => \N__33983\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__6970\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33977\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__33977\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__6968\ : InMux
    port map (
            O => \N__33974\,
            I => \bfn_15_19_0_\
        );

    \I__6967\ : CascadeMux
    port map (
            O => \N__33971\,
            I => \N__33968\
        );

    \I__6966\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33965\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__33965\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__6964\ : InMux
    port map (
            O => \N__33962\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__6963\ : InMux
    port map (
            O => \N__33959\,
            I => \N__33956\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__33956\,
            I => \N__33953\
        );

    \I__6961\ : Span4Mux_h
    port map (
            O => \N__33953\,
            I => \N__33950\
        );

    \I__6960\ : Odrv4
    port map (
            O => \N__33950\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__6959\ : InMux
    port map (
            O => \N__33947\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__6958\ : InMux
    port map (
            O => \N__33944\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__6957\ : InMux
    port map (
            O => \N__33941\,
            I => \N__33938\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__33938\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__6955\ : InMux
    port map (
            O => \N__33935\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__6954\ : InMux
    port map (
            O => \N__33932\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__6953\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33926\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__33926\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__6951\ : InMux
    port map (
            O => \N__33923\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__6950\ : InMux
    port map (
            O => \N__33920\,
            I => \N__33917\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__33917\,
            I => \N__33914\
        );

    \I__6948\ : Odrv4
    port map (
            O => \N__33914\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__6947\ : InMux
    port map (
            O => \N__33911\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__6946\ : InMux
    port map (
            O => \N__33908\,
            I => \N__33905\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__33905\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__6944\ : InMux
    port map (
            O => \N__33902\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__6943\ : InMux
    port map (
            O => \N__33899\,
            I => \N__33896\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__33896\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__6941\ : InMux
    port map (
            O => \N__33893\,
            I => \bfn_15_18_0_\
        );

    \I__6940\ : InMux
    port map (
            O => \N__33890\,
            I => \N__33887\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__33887\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__6938\ : InMux
    port map (
            O => \N__33884\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__6937\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33878\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__33878\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__6935\ : InMux
    port map (
            O => \N__33875\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__6934\ : InMux
    port map (
            O => \N__33872\,
            I => \N__33869\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__33869\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__6932\ : InMux
    port map (
            O => \N__33866\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__6931\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33860\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__33860\,
            I => \N__33857\
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__33857\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__6928\ : InMux
    port map (
            O => \N__33854\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__6927\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33848\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__33848\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__6925\ : InMux
    port map (
            O => \N__33845\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__6924\ : InMux
    port map (
            O => \N__33842\,
            I => \N__33838\
        );

    \I__6923\ : CascadeMux
    port map (
            O => \N__33841\,
            I => \N__33835\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__33838\,
            I => \N__33832\
        );

    \I__6921\ : InMux
    port map (
            O => \N__33835\,
            I => \N__33829\
        );

    \I__6920\ : Span4Mux_h
    port map (
            O => \N__33832\,
            I => \N__33826\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__33829\,
            I => \N__33822\
        );

    \I__6918\ : Span4Mux_v
    port map (
            O => \N__33826\,
            I => \N__33819\
        );

    \I__6917\ : InMux
    port map (
            O => \N__33825\,
            I => \N__33816\
        );

    \I__6916\ : Span4Mux_v
    port map (
            O => \N__33822\,
            I => \N__33813\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__33819\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__33816\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6913\ : Odrv4
    port map (
            O => \N__33813\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6912\ : InMux
    port map (
            O => \N__33806\,
            I => \N__33803\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__33803\,
            I => \N__33800\
        );

    \I__6910\ : Span4Mux_h
    port map (
            O => \N__33800\,
            I => \N__33795\
        );

    \I__6909\ : InMux
    port map (
            O => \N__33799\,
            I => \N__33790\
        );

    \I__6908\ : InMux
    port map (
            O => \N__33798\,
            I => \N__33790\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__33795\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__33790\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__6905\ : InMux
    port map (
            O => \N__33785\,
            I => \N__33782\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__33782\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__6903\ : InMux
    port map (
            O => \N__33779\,
            I => \N__33774\
        );

    \I__6902\ : CascadeMux
    port map (
            O => \N__33778\,
            I => \N__33771\
        );

    \I__6901\ : InMux
    port map (
            O => \N__33777\,
            I => \N__33768\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__33774\,
            I => \N__33765\
        );

    \I__6899\ : InMux
    port map (
            O => \N__33771\,
            I => \N__33762\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__33768\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__6897\ : Odrv4
    port map (
            O => \N__33765\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__33762\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__6895\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33751\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__33754\,
            I => \N__33748\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__33751\,
            I => \N__33745\
        );

    \I__6892\ : InMux
    port map (
            O => \N__33748\,
            I => \N__33742\
        );

    \I__6891\ : Odrv12
    port map (
            O => \N__33745\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__33742\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__6889\ : InMux
    port map (
            O => \N__33737\,
            I => \N__33734\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__33734\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__6887\ : InMux
    port map (
            O => \N__33731\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__6886\ : InMux
    port map (
            O => \N__33728\,
            I => \N__33725\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__33725\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__6884\ : InMux
    port map (
            O => \N__33722\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__6883\ : InMux
    port map (
            O => \N__33719\,
            I => \N__33716\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__33716\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__6881\ : InMux
    port map (
            O => \N__33713\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__6880\ : InMux
    port map (
            O => \N__33710\,
            I => \N__33707\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__33707\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__6878\ : InMux
    port map (
            O => \N__33704\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__6877\ : CascadeMux
    port map (
            O => \N__33701\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_\
        );

    \I__6876\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33695\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__33695\,
            I => \N__33692\
        );

    \I__6874\ : Span4Mux_v
    port map (
            O => \N__33692\,
            I => \N__33687\
        );

    \I__6873\ : InMux
    port map (
            O => \N__33691\,
            I => \N__33684\
        );

    \I__6872\ : InMux
    port map (
            O => \N__33690\,
            I => \N__33681\
        );

    \I__6871\ : Odrv4
    port map (
            O => \N__33687\,
            I => \elapsed_time_ns_1_RNIPFL2M1_0_1\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__33684\,
            I => \elapsed_time_ns_1_RNIPFL2M1_0_1\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__33681\,
            I => \elapsed_time_ns_1_RNIPFL2M1_0_1\
        );

    \I__6868\ : CascadeMux
    port map (
            O => \N__33674\,
            I => \elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_\
        );

    \I__6867\ : InMux
    port map (
            O => \N__33671\,
            I => \N__33668\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__33668\,
            I => \N__33665\
        );

    \I__6865\ : Span4Mux_v
    port map (
            O => \N__33665\,
            I => \N__33661\
        );

    \I__6864\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33658\
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__33661\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_0_1Z0Z_1\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__33658\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_0_1Z0Z_1\
        );

    \I__6861\ : CascadeMux
    port map (
            O => \N__33653\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\
        );

    \I__6860\ : InMux
    port map (
            O => \N__33650\,
            I => \N__33646\
        );

    \I__6859\ : CascadeMux
    port map (
            O => \N__33649\,
            I => \N__33643\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__33646\,
            I => \N__33640\
        );

    \I__6857\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33637\
        );

    \I__6856\ : Span4Mux_h
    port map (
            O => \N__33640\,
            I => \N__33634\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__33637\,
            I => \N__33630\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__33634\,
            I => \N__33627\
        );

    \I__6853\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33624\
        );

    \I__6852\ : Span4Mux_v
    port map (
            O => \N__33630\,
            I => \N__33621\
        );

    \I__6851\ : Odrv4
    port map (
            O => \N__33627\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__33624\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__33621\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6848\ : InMux
    port map (
            O => \N__33614\,
            I => \N__33609\
        );

    \I__6847\ : InMux
    port map (
            O => \N__33613\,
            I => \N__33604\
        );

    \I__6846\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33604\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__33609\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__33604\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6843\ : CascadeMux
    port map (
            O => \N__33599\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_\
        );

    \I__6842\ : InMux
    port map (
            O => \N__33596\,
            I => \N__33593\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__33593\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__6840\ : CascadeMux
    port map (
            O => \N__33590\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\
        );

    \I__6839\ : CascadeMux
    port map (
            O => \N__33587\,
            I => \phase_controller_inst1.stoper_tr.N_251_cascade_\
        );

    \I__6838\ : CascadeMux
    port map (
            O => \N__33584\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5_cascade_\
        );

    \I__6837\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33578\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__33578\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3Z0Z_2\
        );

    \I__6835\ : CascadeMux
    port map (
            O => \N__33575\,
            I => \phase_controller_inst1.stoper_tr.N_241_cascade_\
        );

    \I__6834\ : InMux
    port map (
            O => \N__33572\,
            I => \N__33569\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__33569\,
            I => \N__33566\
        );

    \I__6832\ : Odrv12
    port map (
            O => \N__33566\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\
        );

    \I__6831\ : InMux
    port map (
            O => \N__33563\,
            I => \N__33560\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__33560\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\
        );

    \I__6829\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33554\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__33554\,
            I => \delay_measurement_inst.delay_tr_timer.N_381\
        );

    \I__6827\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33547\
        );

    \I__6826\ : InMux
    port map (
            O => \N__33550\,
            I => \N__33544\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__33547\,
            I => \delay_measurement_inst.delay_tr_timer.N_359_1\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__33544\,
            I => \delay_measurement_inst.delay_tr_timer.N_359_1\
        );

    \I__6823\ : CascadeMux
    port map (
            O => \N__33539\,
            I => \delay_measurement_inst.delay_tr_timer.N_381_cascade_\
        );

    \I__6822\ : CascadeMux
    port map (
            O => \N__33536\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\
        );

    \I__6821\ : CascadeMux
    port map (
            O => \N__33533\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\
        );

    \I__6820\ : CascadeMux
    port map (
            O => \N__33530\,
            I => \N__33527\
        );

    \I__6819\ : InMux
    port map (
            O => \N__33527\,
            I => \N__33523\
        );

    \I__6818\ : InMux
    port map (
            O => \N__33526\,
            I => \N__33520\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__33523\,
            I => \N__33517\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__33520\,
            I => \N__33511\
        );

    \I__6815\ : Span4Mux_v
    port map (
            O => \N__33517\,
            I => \N__33511\
        );

    \I__6814\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33508\
        );

    \I__6813\ : Odrv4
    port map (
            O => \N__33511\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__33508\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__6811\ : InMux
    port map (
            O => \N__33503\,
            I => \N__33500\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__33500\,
            I => \N__33497\
        );

    \I__6809\ : Span4Mux_v
    port map (
            O => \N__33497\,
            I => \N__33494\
        );

    \I__6808\ : Odrv4
    port map (
            O => \N__33494\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\
        );

    \I__6807\ : CascadeMux
    port map (
            O => \N__33491\,
            I => \N__33488\
        );

    \I__6806\ : InMux
    port map (
            O => \N__33488\,
            I => \N__33485\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__33485\,
            I => \N__33482\
        );

    \I__6804\ : Odrv4
    port map (
            O => \N__33482\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__33479\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_\
        );

    \I__6802\ : CascadeMux
    port map (
            O => \N__33476\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\
        );

    \I__6801\ : InMux
    port map (
            O => \N__33473\,
            I => \N__33470\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__33470\,
            I => \elapsed_time_ns_1_RNI3JIF91_0_29\
        );

    \I__6799\ : CascadeMux
    port map (
            O => \N__33467\,
            I => \N__33464\
        );

    \I__6798\ : InMux
    port map (
            O => \N__33464\,
            I => \N__33460\
        );

    \I__6797\ : InMux
    port map (
            O => \N__33463\,
            I => \N__33457\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__33460\,
            I => \elapsed_time_ns_1_RNIRBJF91_0_30\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__33457\,
            I => \elapsed_time_ns_1_RNIRBJF91_0_30\
        );

    \I__6794\ : InMux
    port map (
            O => \N__33452\,
            I => \N__33446\
        );

    \I__6793\ : InMux
    port map (
            O => \N__33451\,
            I => \N__33446\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__33446\,
            I => \elapsed_time_ns_1_RNIRAIF91_0_21\
        );

    \I__6791\ : CascadeMux
    port map (
            O => \N__33443\,
            I => \elapsed_time_ns_1_RNI3JIF91_0_29_cascade_\
        );

    \I__6790\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33436\
        );

    \I__6789\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33433\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__33436\,
            I => \elapsed_time_ns_1_RNIQ9IF91_0_20\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__33433\,
            I => \elapsed_time_ns_1_RNIQ9IF91_0_20\
        );

    \I__6786\ : InMux
    port map (
            O => \N__33428\,
            I => \N__33422\
        );

    \I__6785\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33422\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__33422\,
            I => \N__33419\
        );

    \I__6783\ : Odrv4
    port map (
            O => \N__33419\,
            I => \elapsed_time_ns_1_RNISBIF91_0_22\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__33416\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_o5_7Z0Z_15_cascade_\
        );

    \I__6781\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33410\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__33410\,
            I => \N__33407\
        );

    \I__6779\ : Span4Mux_h
    port map (
            O => \N__33407\,
            I => \N__33404\
        );

    \I__6778\ : Span4Mux_v
    port map (
            O => \N__33404\,
            I => \N__33401\
        );

    \I__6777\ : Odrv4
    port map (
            O => \N__33401\,
            I => \current_shift_inst.PI_CTRL.integrator_i_27\
        );

    \I__6776\ : CascadeMux
    port map (
            O => \N__33398\,
            I => \N__33395\
        );

    \I__6775\ : InMux
    port map (
            O => \N__33395\,
            I => \N__33392\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__33392\,
            I => \N__33389\
        );

    \I__6773\ : Span4Mux_h
    port map (
            O => \N__33389\,
            I => \N__33386\
        );

    \I__6772\ : Span4Mux_v
    port map (
            O => \N__33386\,
            I => \N__33383\
        );

    \I__6771\ : Odrv4
    port map (
            O => \N__33383\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\
        );

    \I__6770\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33377\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__33377\,
            I => \N__33374\
        );

    \I__6768\ : Span4Mux_h
    port map (
            O => \N__33374\,
            I => \N__33371\
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__33371\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__6766\ : InMux
    port map (
            O => \N__33368\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\
        );

    \I__6765\ : CascadeMux
    port map (
            O => \N__33365\,
            I => \N__33362\
        );

    \I__6764\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33359\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__33359\,
            I => \N__33356\
        );

    \I__6762\ : Span12Mux_v
    port map (
            O => \N__33356\,
            I => \N__33353\
        );

    \I__6761\ : Odrv12
    port map (
            O => \N__33353\,
            I => \current_shift_inst.PI_CTRL.integrator_i_28\
        );

    \I__6760\ : InMux
    port map (
            O => \N__33350\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\
        );

    \I__6759\ : CascadeMux
    port map (
            O => \N__33347\,
            I => \N__33344\
        );

    \I__6758\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33341\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__33341\,
            I => \N__33338\
        );

    \I__6756\ : Odrv12
    port map (
            O => \N__33338\,
            I => \current_shift_inst.PI_CTRL.integrator_i_29\
        );

    \I__6755\ : InMux
    port map (
            O => \N__33335\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\
        );

    \I__6754\ : InMux
    port map (
            O => \N__33332\,
            I => \N__33327\
        );

    \I__6753\ : InMux
    port map (
            O => \N__33331\,
            I => \N__33322\
        );

    \I__6752\ : InMux
    port map (
            O => \N__33330\,
            I => \N__33322\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__33327\,
            I => \N__33317\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__33322\,
            I => \N__33317\
        );

    \I__6749\ : Span4Mux_h
    port map (
            O => \N__33317\,
            I => \N__33314\
        );

    \I__6748\ : Odrv4
    port map (
            O => \N__33314\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_0_12\
        );

    \I__6747\ : CascadeMux
    port map (
            O => \N__33311\,
            I => \N__33308\
        );

    \I__6746\ : InMux
    port map (
            O => \N__33308\,
            I => \N__33305\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__33305\,
            I => \N__33302\
        );

    \I__6744\ : Span4Mux_v
    port map (
            O => \N__33302\,
            I => \N__33299\
        );

    \I__6743\ : Span4Mux_v
    port map (
            O => \N__33299\,
            I => \N__33296\
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__33296\,
            I => \current_shift_inst.PI_CTRL.integrator_i_30\
        );

    \I__6741\ : InMux
    port map (
            O => \N__33293\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\
        );

    \I__6740\ : InMux
    port map (
            O => \N__33290\,
            I => \bfn_15_11_0_\
        );

    \I__6739\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33284\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__33284\,
            I => \N__33281\
        );

    \I__6737\ : Odrv4
    port map (
            O => \N__33281\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6\
        );

    \I__6736\ : CascadeMux
    port map (
            O => \N__33278\,
            I => \delay_measurement_inst.delay_tr_timer.N_363_cascade_\
        );

    \I__6735\ : InMux
    port map (
            O => \N__33275\,
            I => \N__33272\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__33272\,
            I => \N__33269\
        );

    \I__6733\ : Span4Mux_v
    port map (
            O => \N__33269\,
            I => \N__33265\
        );

    \I__6732\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33261\
        );

    \I__6731\ : Span4Mux_h
    port map (
            O => \N__33265\,
            I => \N__33258\
        );

    \I__6730\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33255\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__33261\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__6728\ : Odrv4
    port map (
            O => \N__33258\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__33255\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__6726\ : CascadeMux
    port map (
            O => \N__33248\,
            I => \N__33245\
        );

    \I__6725\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33242\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__33242\,
            I => \N__33239\
        );

    \I__6723\ : Span4Mux_h
    port map (
            O => \N__33239\,
            I => \N__33236\
        );

    \I__6722\ : Odrv4
    port map (
            O => \N__33236\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\
        );

    \I__6721\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33230\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__33230\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\
        );

    \I__6719\ : InMux
    port map (
            O => \N__33227\,
            I => \N__33224\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__33224\,
            I => \N__33221\
        );

    \I__6717\ : Odrv4
    port map (
            O => \N__33221\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__6716\ : InMux
    port map (
            O => \N__33218\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\
        );

    \I__6715\ : InMux
    port map (
            O => \N__33215\,
            I => \N__33212\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__33212\,
            I => \N__33209\
        );

    \I__6713\ : Span4Mux_v
    port map (
            O => \N__33209\,
            I => \N__33206\
        );

    \I__6712\ : Span4Mux_v
    port map (
            O => \N__33206\,
            I => \N__33203\
        );

    \I__6711\ : Odrv4
    port map (
            O => \N__33203\,
            I => \current_shift_inst.PI_CTRL.integrator_i_20\
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__33200\,
            I => \N__33197\
        );

    \I__6709\ : InMux
    port map (
            O => \N__33197\,
            I => \N__33194\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__33194\,
            I => \N__33191\
        );

    \I__6707\ : Odrv4
    port map (
            O => \N__33191\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\
        );

    \I__6706\ : CascadeMux
    port map (
            O => \N__33188\,
            I => \N__33185\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33182\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__33182\,
            I => \N__33179\
        );

    \I__6703\ : Odrv12
    port map (
            O => \N__33179\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__6702\ : InMux
    port map (
            O => \N__33176\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\
        );

    \I__6701\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33170\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__33170\,
            I => \N__33167\
        );

    \I__6699\ : Span4Mux_v
    port map (
            O => \N__33167\,
            I => \N__33164\
        );

    \I__6698\ : Odrv4
    port map (
            O => \N__33164\,
            I => \current_shift_inst.PI_CTRL.integrator_i_21\
        );

    \I__6697\ : CascadeMux
    port map (
            O => \N__33161\,
            I => \N__33158\
        );

    \I__6696\ : InMux
    port map (
            O => \N__33158\,
            I => \N__33155\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__33155\,
            I => \N__33152\
        );

    \I__6694\ : Span4Mux_h
    port map (
            O => \N__33152\,
            I => \N__33149\
        );

    \I__6693\ : Odrv4
    port map (
            O => \N__33149\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\
        );

    \I__6692\ : InMux
    port map (
            O => \N__33146\,
            I => \N__33143\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__33143\,
            I => \N__33140\
        );

    \I__6690\ : Odrv12
    port map (
            O => \N__33140\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__6689\ : InMux
    port map (
            O => \N__33137\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\
        );

    \I__6688\ : InMux
    port map (
            O => \N__33134\,
            I => \N__33131\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__33131\,
            I => \N__33128\
        );

    \I__6686\ : Span4Mux_v
    port map (
            O => \N__33128\,
            I => \N__33125\
        );

    \I__6685\ : Odrv4
    port map (
            O => \N__33125\,
            I => \current_shift_inst.PI_CTRL.integrator_i_22\
        );

    \I__6684\ : CascadeMux
    port map (
            O => \N__33122\,
            I => \N__33119\
        );

    \I__6683\ : InMux
    port map (
            O => \N__33119\,
            I => \N__33116\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__33116\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__33113\,
            I => \N__33110\
        );

    \I__6680\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33107\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__33107\,
            I => \N__33104\
        );

    \I__6678\ : Span4Mux_h
    port map (
            O => \N__33104\,
            I => \N__33101\
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__33101\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__6676\ : InMux
    port map (
            O => \N__33098\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\
        );

    \I__6675\ : CascadeMux
    port map (
            O => \N__33095\,
            I => \N__33092\
        );

    \I__6674\ : InMux
    port map (
            O => \N__33092\,
            I => \N__33089\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__33089\,
            I => \current_shift_inst.PI_CTRL.integrator_i_23\
        );

    \I__6672\ : InMux
    port map (
            O => \N__33086\,
            I => \bfn_15_10_0_\
        );

    \I__6671\ : CascadeMux
    port map (
            O => \N__33083\,
            I => \N__33080\
        );

    \I__6670\ : InMux
    port map (
            O => \N__33080\,
            I => \N__33077\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__33077\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\
        );

    \I__6668\ : InMux
    port map (
            O => \N__33074\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\
        );

    \I__6667\ : InMux
    port map (
            O => \N__33071\,
            I => \N__33068\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__33068\,
            I => \N__33065\
        );

    \I__6665\ : Span4Mux_v
    port map (
            O => \N__33065\,
            I => \N__33062\
        );

    \I__6664\ : Odrv4
    port map (
            O => \N__33062\,
            I => \current_shift_inst.PI_CTRL.integrator_i_25\
        );

    \I__6663\ : InMux
    port map (
            O => \N__33059\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\
        );

    \I__6662\ : InMux
    port map (
            O => \N__33056\,
            I => \N__33053\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__33053\,
            I => \current_shift_inst.PI_CTRL.integrator_i_26\
        );

    \I__6660\ : CascadeMux
    port map (
            O => \N__33050\,
            I => \N__33047\
        );

    \I__6659\ : InMux
    port map (
            O => \N__33047\,
            I => \N__33044\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__33044\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\
        );

    \I__6657\ : InMux
    port map (
            O => \N__33041\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\
        );

    \I__6656\ : InMux
    port map (
            O => \N__33038\,
            I => \N__33035\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__33035\,
            I => \N__33032\
        );

    \I__6654\ : Span4Mux_h
    port map (
            O => \N__33032\,
            I => \N__33029\
        );

    \I__6653\ : Odrv4
    port map (
            O => \N__33029\,
            I => \current_shift_inst.PI_CTRL.integrator_i_12\
        );

    \I__6652\ : CascadeMux
    port map (
            O => \N__33026\,
            I => \N__33023\
        );

    \I__6651\ : InMux
    port map (
            O => \N__33023\,
            I => \N__33020\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__33020\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\
        );

    \I__6649\ : InMux
    port map (
            O => \N__33017\,
            I => \N__33014\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__33014\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__6647\ : InMux
    port map (
            O => \N__33011\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\
        );

    \I__6646\ : InMux
    port map (
            O => \N__33008\,
            I => \N__33005\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__33005\,
            I => \N__33002\
        );

    \I__6644\ : Span12Mux_h
    port map (
            O => \N__33002\,
            I => \N__32999\
        );

    \I__6643\ : Odrv12
    port map (
            O => \N__32999\,
            I => \current_shift_inst.PI_CTRL.integrator_i_13\
        );

    \I__6642\ : CascadeMux
    port map (
            O => \N__32996\,
            I => \N__32993\
        );

    \I__6641\ : InMux
    port map (
            O => \N__32993\,
            I => \N__32990\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__32990\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\
        );

    \I__6639\ : CascadeMux
    port map (
            O => \N__32987\,
            I => \N__32984\
        );

    \I__6638\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32981\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__32981\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__6636\ : InMux
    port map (
            O => \N__32978\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\
        );

    \I__6635\ : CascadeMux
    port map (
            O => \N__32975\,
            I => \N__32972\
        );

    \I__6634\ : InMux
    port map (
            O => \N__32972\,
            I => \N__32969\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__32969\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\
        );

    \I__6632\ : CascadeMux
    port map (
            O => \N__32966\,
            I => \N__32963\
        );

    \I__6631\ : InMux
    port map (
            O => \N__32963\,
            I => \N__32960\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__32960\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__6629\ : InMux
    port map (
            O => \N__32957\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\
        );

    \I__6628\ : InMux
    port map (
            O => \N__32954\,
            I => \N__32951\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__32951\,
            I => \current_shift_inst.PI_CTRL.integrator_i_15\
        );

    \I__6626\ : CascadeMux
    port map (
            O => \N__32948\,
            I => \N__32945\
        );

    \I__6625\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32942\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__32942\,
            I => \N__32939\
        );

    \I__6623\ : Odrv12
    port map (
            O => \N__32939\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\
        );

    \I__6622\ : InMux
    port map (
            O => \N__32936\,
            I => \N__32933\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__32933\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__6620\ : InMux
    port map (
            O => \N__32930\,
            I => \bfn_15_9_0_\
        );

    \I__6619\ : InMux
    port map (
            O => \N__32927\,
            I => \N__32924\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__32924\,
            I => \N__32921\
        );

    \I__6617\ : Span4Mux_h
    port map (
            O => \N__32921\,
            I => \N__32918\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__32918\,
            I => \current_shift_inst.PI_CTRL.integrator_i_16\
        );

    \I__6615\ : CascadeMux
    port map (
            O => \N__32915\,
            I => \N__32912\
        );

    \I__6614\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32909\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__32909\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\
        );

    \I__6612\ : InMux
    port map (
            O => \N__32906\,
            I => \N__32903\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__32903\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__6610\ : InMux
    port map (
            O => \N__32900\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\
        );

    \I__6609\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32894\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__32894\,
            I => \N__32891\
        );

    \I__6607\ : Span4Mux_h
    port map (
            O => \N__32891\,
            I => \N__32888\
        );

    \I__6606\ : Odrv4
    port map (
            O => \N__32888\,
            I => \current_shift_inst.PI_CTRL.integrator_i_17\
        );

    \I__6605\ : CascadeMux
    port map (
            O => \N__32885\,
            I => \N__32882\
        );

    \I__6604\ : InMux
    port map (
            O => \N__32882\,
            I => \N__32879\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__32879\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\
        );

    \I__6602\ : InMux
    port map (
            O => \N__32876\,
            I => \N__32873\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__32873\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__6600\ : InMux
    port map (
            O => \N__32870\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\
        );

    \I__6599\ : InMux
    port map (
            O => \N__32867\,
            I => \N__32864\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__32864\,
            I => \N__32861\
        );

    \I__6597\ : Odrv12
    port map (
            O => \N__32861\,
            I => \current_shift_inst.PI_CTRL.integrator_i_18\
        );

    \I__6596\ : CascadeMux
    port map (
            O => \N__32858\,
            I => \N__32855\
        );

    \I__6595\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32852\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__32852\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\
        );

    \I__6593\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32846\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__32846\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__6591\ : InMux
    port map (
            O => \N__32843\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\
        );

    \I__6590\ : InMux
    port map (
            O => \N__32840\,
            I => \N__32837\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__32837\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\
        );

    \I__6588\ : CascadeMux
    port map (
            O => \N__32834\,
            I => \N__32831\
        );

    \I__6587\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32828\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__32828\,
            I => \N__32825\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__32825\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\
        );

    \I__6584\ : CascadeMux
    port map (
            O => \N__32822\,
            I => \N__32819\
        );

    \I__6583\ : InMux
    port map (
            O => \N__32819\,
            I => \N__32816\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__32816\,
            I => \N__32813\
        );

    \I__6581\ : Odrv4
    port map (
            O => \N__32813\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__6580\ : InMux
    port map (
            O => \N__32810\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\
        );

    \I__6579\ : InMux
    port map (
            O => \N__32807\,
            I => \N__32804\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__32804\,
            I => \N__32801\
        );

    \I__6577\ : Span4Mux_h
    port map (
            O => \N__32801\,
            I => \N__32798\
        );

    \I__6576\ : Odrv4
    port map (
            O => \N__32798\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\
        );

    \I__6575\ : CascadeMux
    port map (
            O => \N__32795\,
            I => \N__32792\
        );

    \I__6574\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32789\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__32789\,
            I => \N__32786\
        );

    \I__6572\ : Span12Mux_v
    port map (
            O => \N__32786\,
            I => \N__32783\
        );

    \I__6571\ : Odrv12
    port map (
            O => \N__32783\,
            I => \current_shift_inst.PI_CTRL.integrator_i_5\
        );

    \I__6570\ : InMux
    port map (
            O => \N__32780\,
            I => \N__32777\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__32777\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__6568\ : InMux
    port map (
            O => \N__32774\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\
        );

    \I__6567\ : InMux
    port map (
            O => \N__32771\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\
        );

    \I__6566\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32765\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__32765\,
            I => \current_shift_inst.PI_CTRL.integrator_i_7\
        );

    \I__6564\ : CascadeMux
    port map (
            O => \N__32762\,
            I => \N__32759\
        );

    \I__6563\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32756\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__32756\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\
        );

    \I__6561\ : InMux
    port map (
            O => \N__32753\,
            I => \N__32750\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__32750\,
            I => \N__32747\
        );

    \I__6559\ : Odrv4
    port map (
            O => \N__32747\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__6558\ : InMux
    port map (
            O => \N__32744\,
            I => \bfn_15_8_0_\
        );

    \I__6557\ : InMux
    port map (
            O => \N__32741\,
            I => \N__32738\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__32738\,
            I => \N__32735\
        );

    \I__6555\ : Odrv12
    port map (
            O => \N__32735\,
            I => \current_shift_inst.PI_CTRL.integrator_i_8\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__32732\,
            I => \N__32729\
        );

    \I__6553\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32726\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__32726\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\
        );

    \I__6551\ : CascadeMux
    port map (
            O => \N__32723\,
            I => \N__32720\
        );

    \I__6550\ : InMux
    port map (
            O => \N__32720\,
            I => \N__32717\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__32717\,
            I => \N__32714\
        );

    \I__6548\ : Span4Mux_h
    port map (
            O => \N__32714\,
            I => \N__32711\
        );

    \I__6547\ : Odrv4
    port map (
            O => \N__32711\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__6546\ : InMux
    port map (
            O => \N__32708\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\
        );

    \I__6545\ : InMux
    port map (
            O => \N__32705\,
            I => \N__32702\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__32702\,
            I => \N__32699\
        );

    \I__6543\ : Odrv4
    port map (
            O => \N__32699\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\
        );

    \I__6542\ : CascadeMux
    port map (
            O => \N__32696\,
            I => \N__32693\
        );

    \I__6541\ : InMux
    port map (
            O => \N__32693\,
            I => \N__32690\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__32690\,
            I => \N__32687\
        );

    \I__6539\ : Span12Mux_v
    port map (
            O => \N__32687\,
            I => \N__32684\
        );

    \I__6538\ : Odrv12
    port map (
            O => \N__32684\,
            I => \current_shift_inst.PI_CTRL.integrator_i_9\
        );

    \I__6537\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32678\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__32678\,
            I => \N__32675\
        );

    \I__6535\ : Odrv4
    port map (
            O => \N__32675\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__6534\ : InMux
    port map (
            O => \N__32672\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\
        );

    \I__6533\ : CascadeMux
    port map (
            O => \N__32669\,
            I => \N__32666\
        );

    \I__6532\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32663\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__32663\,
            I => \N__32660\
        );

    \I__6530\ : Span4Mux_h
    port map (
            O => \N__32660\,
            I => \N__32657\
        );

    \I__6529\ : Odrv4
    port map (
            O => \N__32657\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\
        );

    \I__6528\ : InMux
    port map (
            O => \N__32654\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\
        );

    \I__6527\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32648\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__32648\,
            I => \N__32645\
        );

    \I__6525\ : Span4Mux_h
    port map (
            O => \N__32645\,
            I => \N__32642\
        );

    \I__6524\ : Span4Mux_h
    port map (
            O => \N__32642\,
            I => \N__32639\
        );

    \I__6523\ : Odrv4
    port map (
            O => \N__32639\,
            I => \current_shift_inst.PI_CTRL.integrator_i_11\
        );

    \I__6522\ : CascadeMux
    port map (
            O => \N__32636\,
            I => \N__32633\
        );

    \I__6521\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32630\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__32630\,
            I => \N__32627\
        );

    \I__6519\ : Span4Mux_h
    port map (
            O => \N__32627\,
            I => \N__32624\
        );

    \I__6518\ : Odrv4
    port map (
            O => \N__32624\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\
        );

    \I__6517\ : InMux
    port map (
            O => \N__32621\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\
        );

    \I__6516\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32614\
        );

    \I__6515\ : CascadeMux
    port map (
            O => \N__32617\,
            I => \N__32609\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__32614\,
            I => \N__32605\
        );

    \I__6513\ : InMux
    port map (
            O => \N__32613\,
            I => \N__32602\
        );

    \I__6512\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32599\
        );

    \I__6511\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32596\
        );

    \I__6510\ : InMux
    port map (
            O => \N__32608\,
            I => \N__32593\
        );

    \I__6509\ : Span4Mux_h
    port map (
            O => \N__32605\,
            I => \N__32590\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__32602\,
            I => \N__32587\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__32599\,
            I => \N__32582\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__32596\,
            I => \N__32582\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__32593\,
            I => \N__32575\
        );

    \I__6504\ : Span4Mux_h
    port map (
            O => \N__32590\,
            I => \N__32575\
        );

    \I__6503\ : Span4Mux_v
    port map (
            O => \N__32587\,
            I => \N__32575\
        );

    \I__6502\ : Span4Mux_h
    port map (
            O => \N__32582\,
            I => \N__32572\
        );

    \I__6501\ : Span4Mux_v
    port map (
            O => \N__32575\,
            I => \N__32569\
        );

    \I__6500\ : Odrv4
    port map (
            O => \N__32572\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__6499\ : Odrv4
    port map (
            O => \N__32569\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__6498\ : CascadeMux
    port map (
            O => \N__32564\,
            I => \N__32561\
        );

    \I__6497\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32558\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__32558\,
            I => \N__32553\
        );

    \I__6495\ : CascadeMux
    port map (
            O => \N__32557\,
            I => \N__32550\
        );

    \I__6494\ : InMux
    port map (
            O => \N__32556\,
            I => \N__32546\
        );

    \I__6493\ : Span4Mux_h
    port map (
            O => \N__32553\,
            I => \N__32543\
        );

    \I__6492\ : InMux
    port map (
            O => \N__32550\,
            I => \N__32540\
        );

    \I__6491\ : InMux
    port map (
            O => \N__32549\,
            I => \N__32537\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__32546\,
            I => \N__32534\
        );

    \I__6489\ : Span4Mux_v
    port map (
            O => \N__32543\,
            I => \N__32526\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__32540\,
            I => \N__32526\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__32537\,
            I => \N__32526\
        );

    \I__6486\ : Span4Mux_v
    port map (
            O => \N__32534\,
            I => \N__32523\
        );

    \I__6485\ : InMux
    port map (
            O => \N__32533\,
            I => \N__32520\
        );

    \I__6484\ : Span4Mux_h
    port map (
            O => \N__32526\,
            I => \N__32517\
        );

    \I__6483\ : Odrv4
    port map (
            O => \N__32523\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__32520\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__6481\ : Odrv4
    port map (
            O => \N__32517\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__6480\ : InMux
    port map (
            O => \N__32510\,
            I => \N__32504\
        );

    \I__6479\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32501\
        );

    \I__6478\ : InMux
    port map (
            O => \N__32508\,
            I => \N__32498\
        );

    \I__6477\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32495\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__32504\,
            I => \N__32492\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__32501\,
            I => \N__32488\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__32498\,
            I => \N__32483\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__32495\,
            I => \N__32483\
        );

    \I__6472\ : Span12Mux_h
    port map (
            O => \N__32492\,
            I => \N__32480\
        );

    \I__6471\ : InMux
    port map (
            O => \N__32491\,
            I => \N__32477\
        );

    \I__6470\ : Span4Mux_v
    port map (
            O => \N__32488\,
            I => \N__32472\
        );

    \I__6469\ : Span4Mux_h
    port map (
            O => \N__32483\,
            I => \N__32472\
        );

    \I__6468\ : Odrv12
    port map (
            O => \N__32480\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__32477\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__6466\ : Odrv4
    port map (
            O => \N__32472\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__6465\ : CascadeMux
    port map (
            O => \N__32465\,
            I => \N__32462\
        );

    \I__6464\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32458\
        );

    \I__6463\ : InMux
    port map (
            O => \N__32461\,
            I => \N__32455\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__32458\,
            I => \N__32450\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__32455\,
            I => \N__32450\
        );

    \I__6460\ : Span4Mux_h
    port map (
            O => \N__32450\,
            I => \N__32447\
        );

    \I__6459\ : Odrv4
    port map (
            O => \N__32447\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_12\
        );

    \I__6458\ : InMux
    port map (
            O => \N__32444\,
            I => \N__32440\
        );

    \I__6457\ : InMux
    port map (
            O => \N__32443\,
            I => \N__32437\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__32440\,
            I => \N__32434\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__32437\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__6454\ : Odrv4
    port map (
            O => \N__32434\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__6453\ : CascadeMux
    port map (
            O => \N__32429\,
            I => \N__32426\
        );

    \I__6452\ : InMux
    port map (
            O => \N__32426\,
            I => \N__32423\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__32423\,
            I => \N__32420\
        );

    \I__6450\ : Span4Mux_h
    port map (
            O => \N__32420\,
            I => \N__32417\
        );

    \I__6449\ : Odrv4
    port map (
            O => \N__32417\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__32414\,
            I => \N__32411\
        );

    \I__6447\ : InMux
    port map (
            O => \N__32411\,
            I => \N__32408\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__32408\,
            I => \N__32403\
        );

    \I__6445\ : InMux
    port map (
            O => \N__32407\,
            I => \N__32400\
        );

    \I__6444\ : InMux
    port map (
            O => \N__32406\,
            I => \N__32397\
        );

    \I__6443\ : Span4Mux_v
    port map (
            O => \N__32403\,
            I => \N__32394\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__32400\,
            I => \N__32391\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__32397\,
            I => \N__32388\
        );

    \I__6440\ : Span4Mux_h
    port map (
            O => \N__32394\,
            I => \N__32385\
        );

    \I__6439\ : Span4Mux_h
    port map (
            O => \N__32391\,
            I => \N__32380\
        );

    \I__6438\ : Span4Mux_v
    port map (
            O => \N__32388\,
            I => \N__32380\
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__32385\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__6436\ : Odrv4
    port map (
            O => \N__32380\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__6435\ : InMux
    port map (
            O => \N__32375\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\
        );

    \I__6434\ : InMux
    port map (
            O => \N__32372\,
            I => \N__32369\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__32369\,
            I => \N__32366\
        );

    \I__6432\ : Span12Mux_s9_v
    port map (
            O => \N__32366\,
            I => \N__32363\
        );

    \I__6431\ : Odrv12
    port map (
            O => \N__32363\,
            I => \current_shift_inst.PI_CTRL.integrator_i_1\
        );

    \I__6430\ : CascadeMux
    port map (
            O => \N__32360\,
            I => \N__32357\
        );

    \I__6429\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32354\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__32354\,
            I => \N__32351\
        );

    \I__6427\ : Span4Mux_h
    port map (
            O => \N__32351\,
            I => \N__32348\
        );

    \I__6426\ : Odrv4
    port map (
            O => \N__32348\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\
        );

    \I__6425\ : CascadeMux
    port map (
            O => \N__32345\,
            I => \N__32342\
        );

    \I__6424\ : InMux
    port map (
            O => \N__32342\,
            I => \N__32339\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__32339\,
            I => \N__32333\
        );

    \I__6422\ : InMux
    port map (
            O => \N__32338\,
            I => \N__32328\
        );

    \I__6421\ : InMux
    port map (
            O => \N__32337\,
            I => \N__32328\
        );

    \I__6420\ : CascadeMux
    port map (
            O => \N__32336\,
            I => \N__32325\
        );

    \I__6419\ : Span4Mux_v
    port map (
            O => \N__32333\,
            I => \N__32322\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__32328\,
            I => \N__32319\
        );

    \I__6417\ : InMux
    port map (
            O => \N__32325\,
            I => \N__32316\
        );

    \I__6416\ : Span4Mux_h
    port map (
            O => \N__32322\,
            I => \N__32311\
        );

    \I__6415\ : Span4Mux_v
    port map (
            O => \N__32319\,
            I => \N__32311\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__32316\,
            I => \N__32308\
        );

    \I__6413\ : Span4Mux_h
    port map (
            O => \N__32311\,
            I => \N__32305\
        );

    \I__6412\ : Odrv12
    port map (
            O => \N__32308\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__6411\ : Odrv4
    port map (
            O => \N__32305\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__6410\ : InMux
    port map (
            O => \N__32300\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\
        );

    \I__6409\ : InMux
    port map (
            O => \N__32297\,
            I => \N__32294\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__32294\,
            I => \N__32291\
        );

    \I__6407\ : Span4Mux_h
    port map (
            O => \N__32291\,
            I => \N__32288\
        );

    \I__6406\ : Odrv4
    port map (
            O => \N__32288\,
            I => \current_shift_inst.PI_CTRL.integrator_i_2\
        );

    \I__6405\ : InMux
    port map (
            O => \N__32285\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\
        );

    \I__6404\ : InMux
    port map (
            O => \N__32282\,
            I => \N__32279\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__32279\,
            I => \N__32276\
        );

    \I__6402\ : Span4Mux_h
    port map (
            O => \N__32276\,
            I => \N__32273\
        );

    \I__6401\ : Odrv4
    port map (
            O => \N__32273\,
            I => \current_shift_inst.PI_CTRL.integrator_i_3\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__32270\,
            I => \N__32267\
        );

    \I__6399\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32264\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__32264\,
            I => \N__32261\
        );

    \I__6397\ : Span4Mux_h
    port map (
            O => \N__32261\,
            I => \N__32258\
        );

    \I__6396\ : Odrv4
    port map (
            O => \N__32258\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\
        );

    \I__6395\ : CascadeMux
    port map (
            O => \N__32255\,
            I => \N__32252\
        );

    \I__6394\ : InMux
    port map (
            O => \N__32252\,
            I => \N__32248\
        );

    \I__6393\ : InMux
    port map (
            O => \N__32251\,
            I => \N__32242\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__32248\,
            I => \N__32239\
        );

    \I__6391\ : InMux
    port map (
            O => \N__32247\,
            I => \N__32236\
        );

    \I__6390\ : InMux
    port map (
            O => \N__32246\,
            I => \N__32233\
        );

    \I__6389\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32230\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__32242\,
            I => \N__32225\
        );

    \I__6387\ : Span4Mux_h
    port map (
            O => \N__32239\,
            I => \N__32225\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__32236\,
            I => \N__32220\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__32233\,
            I => \N__32220\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__32230\,
            I => \N__32217\
        );

    \I__6383\ : Span4Mux_h
    port map (
            O => \N__32225\,
            I => \N__32214\
        );

    \I__6382\ : Span4Mux_h
    port map (
            O => \N__32220\,
            I => \N__32211\
        );

    \I__6381\ : Odrv12
    port map (
            O => \N__32217\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__6380\ : Odrv4
    port map (
            O => \N__32214\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__6379\ : Odrv4
    port map (
            O => \N__32211\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__6378\ : InMux
    port map (
            O => \N__32204\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\
        );

    \I__6377\ : InMux
    port map (
            O => \N__32201\,
            I => \N__32198\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__32198\,
            I => \N__32195\
        );

    \I__6375\ : Odrv12
    port map (
            O => \N__32195\,
            I => \current_shift_inst.PI_CTRL.integrator_i_4\
        );

    \I__6374\ : CascadeMux
    port map (
            O => \N__32192\,
            I => \N__32189\
        );

    \I__6373\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32186\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__32186\,
            I => \N__32183\
        );

    \I__6371\ : Odrv12
    port map (
            O => \N__32183\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__6370\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32171\
        );

    \I__6369\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32171\
        );

    \I__6368\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32171\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__32171\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__6366\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32165\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__32165\,
            I => \N__32162\
        );

    \I__6364\ : Odrv12
    port map (
            O => \N__32162\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3\
        );

    \I__6363\ : CascadeMux
    port map (
            O => \N__32159\,
            I => \N__32156\
        );

    \I__6362\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32153\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__32153\,
            I => \N__32150\
        );

    \I__6360\ : Span4Mux_v
    port map (
            O => \N__32150\,
            I => \N__32147\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__32147\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__6358\ : InMux
    port map (
            O => \N__32144\,
            I => \N__32141\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__32141\,
            I => \N__32138\
        );

    \I__6356\ : Odrv4
    port map (
            O => \N__32138\,
            I => \current_shift_inst.un38_control_input_cry_5_c_RNOZ0\
        );

    \I__6355\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32132\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__32132\,
            I => \N__32129\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__32129\,
            I => \current_shift_inst.un38_control_input_cry_13_c_RNOZ0\
        );

    \I__6352\ : CascadeMux
    port map (
            O => \N__32126\,
            I => \N__32123\
        );

    \I__6351\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32120\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__32120\,
            I => \N__32117\
        );

    \I__6349\ : Span12Mux_h
    port map (
            O => \N__32117\,
            I => \N__32114\
        );

    \I__6348\ : Odrv12
    port map (
            O => \N__32114\,
            I => \current_shift_inst.un38_control_input_cry_8_c_RNOZ0\
        );

    \I__6347\ : CascadeMux
    port map (
            O => \N__32111\,
            I => \N__32108\
        );

    \I__6346\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32105\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__32105\,
            I => \N__32102\
        );

    \I__6344\ : Span4Mux_v
    port map (
            O => \N__32102\,
            I => \N__32099\
        );

    \I__6343\ : Odrv4
    port map (
            O => \N__32099\,
            I => \current_shift_inst.un38_control_input_cry_10_c_RNOZ0\
        );

    \I__6342\ : CascadeMux
    port map (
            O => \N__32096\,
            I => \N__32093\
        );

    \I__6341\ : InMux
    port map (
            O => \N__32093\,
            I => \N__32090\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__32090\,
            I => \N__32087\
        );

    \I__6339\ : Span4Mux_h
    port map (
            O => \N__32087\,
            I => \N__32084\
        );

    \I__6338\ : Odrv4
    port map (
            O => \N__32084\,
            I => \current_shift_inst.un38_control_input_cry_12_c_RNOZ0\
        );

    \I__6337\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32078\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__32078\,
            I => \N__32075\
        );

    \I__6335\ : Span4Mux_h
    port map (
            O => \N__32075\,
            I => \N__32072\
        );

    \I__6334\ : Odrv4
    port map (
            O => \N__32072\,
            I => \current_shift_inst.un38_control_input_cry_15_c_RNOZ0\
        );

    \I__6333\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32066\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__32066\,
            I => \N__32063\
        );

    \I__6331\ : Span4Mux_h
    port map (
            O => \N__32063\,
            I => \N__32060\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__32060\,
            I => \current_shift_inst.un38_control_input_cry_2_c_RNOZ0\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__32057\,
            I => \N__32051\
        );

    \I__6328\ : InMux
    port map (
            O => \N__32056\,
            I => \N__32043\
        );

    \I__6327\ : InMux
    port map (
            O => \N__32055\,
            I => \N__32043\
        );

    \I__6326\ : InMux
    port map (
            O => \N__32054\,
            I => \N__32043\
        );

    \I__6325\ : InMux
    port map (
            O => \N__32051\,
            I => \N__32038\
        );

    \I__6324\ : InMux
    port map (
            O => \N__32050\,
            I => \N__32038\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__32043\,
            I => \N__32035\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__32038\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6321\ : Odrv4
    port map (
            O => \N__32035\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6320\ : CascadeMux
    port map (
            O => \N__32030\,
            I => \N__32026\
        );

    \I__6319\ : InMux
    port map (
            O => \N__32029\,
            I => \N__32016\
        );

    \I__6318\ : InMux
    port map (
            O => \N__32026\,
            I => \N__32016\
        );

    \I__6317\ : InMux
    port map (
            O => \N__32025\,
            I => \N__32016\
        );

    \I__6316\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32011\
        );

    \I__6315\ : InMux
    port map (
            O => \N__32023\,
            I => \N__32011\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__32016\,
            I => \N__32008\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__32011\,
            I => \N__32004\
        );

    \I__6312\ : Span4Mux_h
    port map (
            O => \N__32008\,
            I => \N__32001\
        );

    \I__6311\ : InMux
    port map (
            O => \N__32007\,
            I => \N__31998\
        );

    \I__6310\ : Span4Mux_v
    port map (
            O => \N__32004\,
            I => \N__31995\
        );

    \I__6309\ : Span4Mux_v
    port map (
            O => \N__32001\,
            I => \N__31992\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__31998\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6307\ : Odrv4
    port map (
            O => \N__31995\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__31992\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6305\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31982\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__31982\,
            I => \N__31979\
        );

    \I__6303\ : Span4Mux_v
    port map (
            O => \N__31979\,
            I => \N__31976\
        );

    \I__6302\ : Span4Mux_h
    port map (
            O => \N__31976\,
            I => \N__31973\
        );

    \I__6301\ : Odrv4
    port map (
            O => \N__31973\,
            I => \phase_controller_inst2.stoper_hc.N_45\
        );

    \I__6300\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31967\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__31967\,
            I => \N__31964\
        );

    \I__6298\ : Odrv4
    port map (
            O => \N__31964\,
            I => \phase_controller_inst1.stoper_tr.N_219\
        );

    \I__6297\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31958\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__31958\,
            I => \N__31953\
        );

    \I__6295\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31950\
        );

    \I__6294\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31947\
        );

    \I__6293\ : Span4Mux_v
    port map (
            O => \N__31953\,
            I => \N__31942\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__31950\,
            I => \N__31942\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__31947\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__6290\ : Odrv4
    port map (
            O => \N__31942\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__6289\ : InMux
    port map (
            O => \N__31937\,
            I => \N__31933\
        );

    \I__6288\ : InMux
    port map (
            O => \N__31936\,
            I => \N__31930\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__31933\,
            I => \N__31926\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__31930\,
            I => \N__31923\
        );

    \I__6285\ : InMux
    port map (
            O => \N__31929\,
            I => \N__31920\
        );

    \I__6284\ : Span4Mux_v
    port map (
            O => \N__31926\,
            I => \N__31915\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__31923\,
            I => \N__31915\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__31920\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__6281\ : Odrv4
    port map (
            O => \N__31915\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__6280\ : CascadeMux
    port map (
            O => \N__31910\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__6279\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31904\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__31904\,
            I => \N__31901\
        );

    \I__6277\ : Span4Mux_h
    port map (
            O => \N__31901\,
            I => \N__31898\
        );

    \I__6276\ : Odrv4
    port map (
            O => \N__31898\,
            I => \current_shift_inst.un38_control_input_cry_0_c_RNOZ0\
        );

    \I__6275\ : InMux
    port map (
            O => \N__31895\,
            I => \N__31892\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__31892\,
            I => \N__31889\
        );

    \I__6273\ : Span4Mux_h
    port map (
            O => \N__31889\,
            I => \N__31886\
        );

    \I__6272\ : Odrv4
    port map (
            O => \N__31886\,
            I => \current_shift_inst.un38_control_input_cry_6_c_RNOZ0\
        );

    \I__6271\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31880\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__31880\,
            I => \N__31877\
        );

    \I__6269\ : Span4Mux_h
    port map (
            O => \N__31877\,
            I => \N__31874\
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__31874\,
            I => \current_shift_inst.un38_control_input_cry_9_c_RNOZ0\
        );

    \I__6267\ : CascadeMux
    port map (
            O => \N__31871\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7_cascade_\
        );

    \I__6266\ : CascadeMux
    port map (
            O => \N__31868\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2_cascade_\
        );

    \I__6265\ : InMux
    port map (
            O => \N__31865\,
            I => \N__31860\
        );

    \I__6264\ : CascadeMux
    port map (
            O => \N__31864\,
            I => \N__31851\
        );

    \I__6263\ : CascadeMux
    port map (
            O => \N__31863\,
            I => \N__31848\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__31860\,
            I => \N__31844\
        );

    \I__6261\ : InMux
    port map (
            O => \N__31859\,
            I => \N__31839\
        );

    \I__6260\ : InMux
    port map (
            O => \N__31858\,
            I => \N__31839\
        );

    \I__6259\ : InMux
    port map (
            O => \N__31857\,
            I => \N__31836\
        );

    \I__6258\ : InMux
    port map (
            O => \N__31856\,
            I => \N__31830\
        );

    \I__6257\ : InMux
    port map (
            O => \N__31855\,
            I => \N__31830\
        );

    \I__6256\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31827\
        );

    \I__6255\ : InMux
    port map (
            O => \N__31851\,
            I => \N__31820\
        );

    \I__6254\ : InMux
    port map (
            O => \N__31848\,
            I => \N__31820\
        );

    \I__6253\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31820\
        );

    \I__6252\ : Span4Mux_v
    port map (
            O => \N__31844\,
            I => \N__31813\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__31839\,
            I => \N__31810\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__31836\,
            I => \N__31805\
        );

    \I__6249\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31796\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__31830\,
            I => \N__31793\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__31827\,
            I => \N__31788\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__31820\,
            I => \N__31788\
        );

    \I__6245\ : InMux
    port map (
            O => \N__31819\,
            I => \N__31779\
        );

    \I__6244\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31779\
        );

    \I__6243\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31779\
        );

    \I__6242\ : InMux
    port map (
            O => \N__31816\,
            I => \N__31779\
        );

    \I__6241\ : Sp12to4
    port map (
            O => \N__31813\,
            I => \N__31768\
        );

    \I__6240\ : Span4Mux_h
    port map (
            O => \N__31810\,
            I => \N__31765\
        );

    \I__6239\ : InMux
    port map (
            O => \N__31809\,
            I => \N__31762\
        );

    \I__6238\ : InMux
    port map (
            O => \N__31808\,
            I => \N__31759\
        );

    \I__6237\ : Span12Mux_v
    port map (
            O => \N__31805\,
            I => \N__31756\
        );

    \I__6236\ : InMux
    port map (
            O => \N__31804\,
            I => \N__31747\
        );

    \I__6235\ : InMux
    port map (
            O => \N__31803\,
            I => \N__31747\
        );

    \I__6234\ : InMux
    port map (
            O => \N__31802\,
            I => \N__31747\
        );

    \I__6233\ : InMux
    port map (
            O => \N__31801\,
            I => \N__31747\
        );

    \I__6232\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31742\
        );

    \I__6231\ : InMux
    port map (
            O => \N__31799\,
            I => \N__31742\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__31796\,
            I => \N__31735\
        );

    \I__6229\ : Span4Mux_v
    port map (
            O => \N__31793\,
            I => \N__31735\
        );

    \I__6228\ : Span4Mux_v
    port map (
            O => \N__31788\,
            I => \N__31735\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__31779\,
            I => \N__31732\
        );

    \I__6226\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31723\
        );

    \I__6225\ : InMux
    port map (
            O => \N__31777\,
            I => \N__31723\
        );

    \I__6224\ : InMux
    port map (
            O => \N__31776\,
            I => \N__31723\
        );

    \I__6223\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31723\
        );

    \I__6222\ : InMux
    port map (
            O => \N__31774\,
            I => \N__31714\
        );

    \I__6221\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31714\
        );

    \I__6220\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31714\
        );

    \I__6219\ : InMux
    port map (
            O => \N__31771\,
            I => \N__31714\
        );

    \I__6218\ : Odrv12
    port map (
            O => \N__31768\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6217\ : Odrv4
    port map (
            O => \N__31765\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__31762\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__31759\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6214\ : Odrv12
    port map (
            O => \N__31756\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__31747\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__31742\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__31735\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6210\ : Odrv4
    port map (
            O => \N__31732\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__31723\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__31714\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__6207\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31688\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__31688\,
            I => \N__31684\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__31687\,
            I => \N__31680\
        );

    \I__6204\ : Span4Mux_h
    port map (
            O => \N__31684\,
            I => \N__31676\
        );

    \I__6203\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31673\
        );

    \I__6202\ : InMux
    port map (
            O => \N__31680\,
            I => \N__31670\
        );

    \I__6201\ : InMux
    port map (
            O => \N__31679\,
            I => \N__31667\
        );

    \I__6200\ : Odrv4
    port map (
            O => \N__31676\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__31673\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__31670\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__31667\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6\
        );

    \I__6196\ : CascadeMux
    port map (
            O => \N__31658\,
            I => \N__31654\
        );

    \I__6195\ : CascadeMux
    port map (
            O => \N__31657\,
            I => \N__31651\
        );

    \I__6194\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31646\
        );

    \I__6193\ : InMux
    port map (
            O => \N__31651\,
            I => \N__31642\
        );

    \I__6192\ : CascadeMux
    port map (
            O => \N__31650\,
            I => \N__31639\
        );

    \I__6191\ : CascadeMux
    port map (
            O => \N__31649\,
            I => \N__31634\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__31646\,
            I => \N__31631\
        );

    \I__6189\ : InMux
    port map (
            O => \N__31645\,
            I => \N__31628\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__31642\,
            I => \N__31625\
        );

    \I__6187\ : InMux
    port map (
            O => \N__31639\,
            I => \N__31622\
        );

    \I__6186\ : InMux
    port map (
            O => \N__31638\,
            I => \N__31614\
        );

    \I__6185\ : InMux
    port map (
            O => \N__31637\,
            I => \N__31614\
        );

    \I__6184\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31614\
        );

    \I__6183\ : Sp12to4
    port map (
            O => \N__31631\,
            I => \N__31609\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__31628\,
            I => \N__31609\
        );

    \I__6181\ : Span4Mux_h
    port map (
            O => \N__31625\,
            I => \N__31603\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__31622\,
            I => \N__31603\
        );

    \I__6179\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31600\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__31614\,
            I => \N__31597\
        );

    \I__6177\ : Span12Mux_v
    port map (
            O => \N__31609\,
            I => \N__31594\
        );

    \I__6176\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31591\
        );

    \I__6175\ : Span4Mux_h
    port map (
            O => \N__31603\,
            I => \N__31584\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__31600\,
            I => \N__31584\
        );

    \I__6173\ : Span4Mux_h
    port map (
            O => \N__31597\,
            I => \N__31584\
        );

    \I__6172\ : Odrv12
    port map (
            O => \N__31594\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__31591\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__31584\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__6169\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31574\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__31574\,
            I => \N__31571\
        );

    \I__6167\ : Span4Mux_h
    port map (
            O => \N__31571\,
            I => \N__31567\
        );

    \I__6166\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31563\
        );

    \I__6165\ : Span4Mux_v
    port map (
            O => \N__31567\,
            I => \N__31560\
        );

    \I__6164\ : InMux
    port map (
            O => \N__31566\,
            I => \N__31557\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__31563\,
            I => \N__31554\
        );

    \I__6162\ : Odrv4
    port map (
            O => \N__31560\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__31557\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\
        );

    \I__6160\ : Odrv4
    port map (
            O => \N__31554\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\
        );

    \I__6159\ : InMux
    port map (
            O => \N__31547\,
            I => \N__31544\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__31544\,
            I => \N__31541\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__31541\,
            I => \N__31538\
        );

    \I__6156\ : Odrv4
    port map (
            O => \N__31538\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6\
        );

    \I__6155\ : CascadeMux
    port map (
            O => \N__31535\,
            I => \phase_controller_inst1.stoper_tr.N_235_cascade_\
        );

    \I__6154\ : CascadeMux
    port map (
            O => \N__31532\,
            I => \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3_cascade_\
        );

    \I__6153\ : CEMux
    port map (
            O => \N__31529\,
            I => \N__31523\
        );

    \I__6152\ : CEMux
    port map (
            O => \N__31528\,
            I => \N__31519\
        );

    \I__6151\ : CEMux
    port map (
            O => \N__31527\,
            I => \N__31516\
        );

    \I__6150\ : CEMux
    port map (
            O => \N__31526\,
            I => \N__31513\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__31523\,
            I => \N__31510\
        );

    \I__6148\ : CEMux
    port map (
            O => \N__31522\,
            I => \N__31507\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__31519\,
            I => \N__31504\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__31516\,
            I => \N__31501\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__31513\,
            I => \N__31498\
        );

    \I__6144\ : Span4Mux_v
    port map (
            O => \N__31510\,
            I => \N__31493\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__31507\,
            I => \N__31493\
        );

    \I__6142\ : Span4Mux_h
    port map (
            O => \N__31504\,
            I => \N__31488\
        );

    \I__6141\ : Span4Mux_h
    port map (
            O => \N__31501\,
            I => \N__31488\
        );

    \I__6140\ : Span4Mux_h
    port map (
            O => \N__31498\,
            I => \N__31483\
        );

    \I__6139\ : Span4Mux_h
    port map (
            O => \N__31493\,
            I => \N__31483\
        );

    \I__6138\ : Span4Mux_h
    port map (
            O => \N__31488\,
            I => \N__31480\
        );

    \I__6137\ : Span4Mux_h
    port map (
            O => \N__31483\,
            I => \N__31477\
        );

    \I__6136\ : Odrv4
    port map (
            O => \N__31480\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa_0\
        );

    \I__6135\ : Odrv4
    port map (
            O => \N__31477\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa_0\
        );

    \I__6134\ : InMux
    port map (
            O => \N__31472\,
            I => \N__31467\
        );

    \I__6133\ : CascadeMux
    port map (
            O => \N__31471\,
            I => \N__31464\
        );

    \I__6132\ : InMux
    port map (
            O => \N__31470\,
            I => \N__31459\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__31467\,
            I => \N__31453\
        );

    \I__6130\ : InMux
    port map (
            O => \N__31464\,
            I => \N__31448\
        );

    \I__6129\ : InMux
    port map (
            O => \N__31463\,
            I => \N__31448\
        );

    \I__6128\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31445\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__31459\,
            I => \N__31442\
        );

    \I__6126\ : InMux
    port map (
            O => \N__31458\,
            I => \N__31439\
        );

    \I__6125\ : InMux
    port map (
            O => \N__31457\,
            I => \N__31434\
        );

    \I__6124\ : InMux
    port map (
            O => \N__31456\,
            I => \N__31434\
        );

    \I__6123\ : Span4Mux_v
    port map (
            O => \N__31453\,
            I => \N__31431\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__31448\,
            I => \N__31428\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__31445\,
            I => \N__31423\
        );

    \I__6120\ : Span4Mux_h
    port map (
            O => \N__31442\,
            I => \N__31423\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__31439\,
            I => \N__31420\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__31434\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6117\ : Odrv4
    port map (
            O => \N__31431\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__31428\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6115\ : Odrv4
    port map (
            O => \N__31423\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6114\ : Odrv4
    port map (
            O => \N__31420\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6113\ : SRMux
    port map (
            O => \N__31409\,
            I => \N__31404\
        );

    \I__6112\ : SRMux
    port map (
            O => \N__31408\,
            I => \N__31401\
        );

    \I__6111\ : SRMux
    port map (
            O => \N__31407\,
            I => \N__31397\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__31404\,
            I => \N__31394\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31391\
        );

    \I__6108\ : SRMux
    port map (
            O => \N__31400\,
            I => \N__31388\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__31397\,
            I => \N__31385\
        );

    \I__6106\ : Span4Mux_v
    port map (
            O => \N__31394\,
            I => \N__31378\
        );

    \I__6105\ : Span4Mux_v
    port map (
            O => \N__31391\,
            I => \N__31378\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__31388\,
            I => \N__31378\
        );

    \I__6103\ : Span4Mux_h
    port map (
            O => \N__31385\,
            I => \N__31375\
        );

    \I__6102\ : Sp12to4
    port map (
            O => \N__31378\,
            I => \N__31372\
        );

    \I__6101\ : Span4Mux_h
    port map (
            O => \N__31375\,
            I => \N__31369\
        );

    \I__6100\ : Odrv12
    port map (
            O => \N__31372\,
            I => \phase_controller_inst2.stoper_hc.un1_stoper_state12_1_0_i\
        );

    \I__6099\ : Odrv4
    port map (
            O => \N__31369\,
            I => \phase_controller_inst2.stoper_hc.un1_stoper_state12_1_0_i\
        );

    \I__6098\ : CascadeMux
    port map (
            O => \N__31364\,
            I => \delay_measurement_inst.delay_tr_timer.N_358_cascade_\
        );

    \I__6097\ : CascadeMux
    port map (
            O => \N__31361\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__31358\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9_cascade_\
        );

    \I__6095\ : InMux
    port map (
            O => \N__31355\,
            I => \N__31352\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__31352\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\
        );

    \I__6093\ : InMux
    port map (
            O => \N__31349\,
            I => \N__31345\
        );

    \I__6092\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31342\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__31345\,
            I => \N__31338\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__31342\,
            I => \N__31335\
        );

    \I__6089\ : InMux
    port map (
            O => \N__31341\,
            I => \N__31332\
        );

    \I__6088\ : Span4Mux_h
    port map (
            O => \N__31338\,
            I => \N__31329\
        );

    \I__6087\ : Span4Mux_v
    port map (
            O => \N__31335\,
            I => \N__31326\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__31332\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__6085\ : Odrv4
    port map (
            O => \N__31329\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__6084\ : Odrv4
    port map (
            O => \N__31326\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__6083\ : InMux
    port map (
            O => \N__31319\,
            I => \N__31316\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__31316\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\
        );

    \I__6081\ : CascadeMux
    port map (
            O => \N__31313\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_\
        );

    \I__6080\ : CascadeMux
    port map (
            O => \N__31310\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\
        );

    \I__6079\ : CascadeMux
    port map (
            O => \N__31307\,
            I => \N__31304\
        );

    \I__6078\ : InMux
    port map (
            O => \N__31304\,
            I => \N__31300\
        );

    \I__6077\ : InMux
    port map (
            O => \N__31303\,
            I => \N__31297\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__31300\,
            I => \N__31294\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__31297\,
            I => \N__31288\
        );

    \I__6074\ : Span4Mux_v
    port map (
            O => \N__31294\,
            I => \N__31288\
        );

    \I__6073\ : InMux
    port map (
            O => \N__31293\,
            I => \N__31285\
        );

    \I__6072\ : Odrv4
    port map (
            O => \N__31288\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__31285\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__6070\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31277\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__31277\,
            I => \N__31274\
        );

    \I__6068\ : Span4Mux_v
    port map (
            O => \N__31274\,
            I => \N__31271\
        );

    \I__6067\ : Odrv4
    port map (
            O => \N__31271\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\
        );

    \I__6066\ : InMux
    port map (
            O => \N__31268\,
            I => \N__31264\
        );

    \I__6065\ : InMux
    port map (
            O => \N__31267\,
            I => \N__31260\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__31264\,
            I => \N__31257\
        );

    \I__6063\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31254\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__31260\,
            I => \N__31250\
        );

    \I__6061\ : Span4Mux_h
    port map (
            O => \N__31257\,
            I => \N__31245\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31245\
        );

    \I__6059\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31242\
        );

    \I__6058\ : Span4Mux_v
    port map (
            O => \N__31250\,
            I => \N__31234\
        );

    \I__6057\ : Span4Mux_v
    port map (
            O => \N__31245\,
            I => \N__31234\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__31242\,
            I => \N__31234\
        );

    \I__6055\ : InMux
    port map (
            O => \N__31241\,
            I => \N__31231\
        );

    \I__6054\ : Odrv4
    port map (
            O => \N__31234\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__31231\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__6052\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31222\
        );

    \I__6051\ : InMux
    port map (
            O => \N__31225\,
            I => \N__31219\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__31222\,
            I => \N__31216\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__31219\,
            I => \N__31213\
        );

    \I__6048\ : Span4Mux_v
    port map (
            O => \N__31216\,
            I => \N__31209\
        );

    \I__6047\ : Span4Mux_h
    port map (
            O => \N__31213\,
            I => \N__31206\
        );

    \I__6046\ : InMux
    port map (
            O => \N__31212\,
            I => \N__31203\
        );

    \I__6045\ : Odrv4
    port map (
            O => \N__31209\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6044\ : Odrv4
    port map (
            O => \N__31206\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__31203\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6042\ : InMux
    port map (
            O => \N__31196\,
            I => \N__31193\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__31193\,
            I => \N__31190\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__31190\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_9\
        );

    \I__6039\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31182\
        );

    \I__6038\ : InMux
    port map (
            O => \N__31186\,
            I => \N__31179\
        );

    \I__6037\ : InMux
    port map (
            O => \N__31185\,
            I => \N__31176\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__31182\,
            I => \N__31173\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__31179\,
            I => \N__31170\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__31176\,
            I => \N__31163\
        );

    \I__6033\ : Span4Mux_v
    port map (
            O => \N__31173\,
            I => \N__31163\
        );

    \I__6032\ : Span4Mux_v
    port map (
            O => \N__31170\,
            I => \N__31163\
        );

    \I__6031\ : Odrv4
    port map (
            O => \N__31163\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__6030\ : InMux
    port map (
            O => \N__31160\,
            I => \N__31157\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__31157\,
            I => \N__31154\
        );

    \I__6028\ : Span4Mux_h
    port map (
            O => \N__31154\,
            I => \N__31151\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__31151\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\
        );

    \I__6026\ : CascadeMux
    port map (
            O => \N__31148\,
            I => \N__31145\
        );

    \I__6025\ : InMux
    port map (
            O => \N__31145\,
            I => \N__31142\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__31142\,
            I => \N__31138\
        );

    \I__6023\ : InMux
    port map (
            O => \N__31141\,
            I => \N__31134\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__31138\,
            I => \N__31131\
        );

    \I__6021\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31128\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__31134\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__6019\ : Odrv4
    port map (
            O => \N__31131\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__31128\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__6017\ : InMux
    port map (
            O => \N__31121\,
            I => \N__31118\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__31118\,
            I => \N__31115\
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__31115\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\
        );

    \I__6014\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31108\
        );

    \I__6013\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31105\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__31108\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__31105\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__31100\,
            I => \N__31097\
        );

    \I__6009\ : InMux
    port map (
            O => \N__31097\,
            I => \N__31092\
        );

    \I__6008\ : CascadeMux
    port map (
            O => \N__31096\,
            I => \N__31089\
        );

    \I__6007\ : InMux
    port map (
            O => \N__31095\,
            I => \N__31086\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__31092\,
            I => \N__31082\
        );

    \I__6005\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31079\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__31086\,
            I => \N__31076\
        );

    \I__6003\ : InMux
    port map (
            O => \N__31085\,
            I => \N__31073\
        );

    \I__6002\ : Span4Mux_h
    port map (
            O => \N__31082\,
            I => \N__31070\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__31079\,
            I => \N__31067\
        );

    \I__6000\ : Span4Mux_v
    port map (
            O => \N__31076\,
            I => \N__31060\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__31073\,
            I => \N__31060\
        );

    \I__5998\ : Span4Mux_v
    port map (
            O => \N__31070\,
            I => \N__31060\
        );

    \I__5997\ : Span4Mux_v
    port map (
            O => \N__31067\,
            I => \N__31056\
        );

    \I__5996\ : Span4Mux_h
    port map (
            O => \N__31060\,
            I => \N__31053\
        );

    \I__5995\ : InMux
    port map (
            O => \N__31059\,
            I => \N__31050\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__31056\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__5993\ : Odrv4
    port map (
            O => \N__31053\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__31050\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__31043\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13_cascade_\
        );

    \I__5990\ : InMux
    port map (
            O => \N__31040\,
            I => \N__31037\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__31037\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\
        );

    \I__5988\ : InMux
    port map (
            O => \N__31034\,
            I => \N__31030\
        );

    \I__5987\ : InMux
    port map (
            O => \N__31033\,
            I => \N__31027\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__31030\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__31027\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__5984\ : CascadeMux
    port map (
            O => \N__31022\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14_cascade_\
        );

    \I__5983\ : InMux
    port map (
            O => \N__31019\,
            I => \N__31016\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__31016\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__31013\,
            I => \N__31010\
        );

    \I__5980\ : InMux
    port map (
            O => \N__31010\,
            I => \N__31006\
        );

    \I__5979\ : CascadeMux
    port map (
            O => \N__31009\,
            I => \N__31003\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__31006\,
            I => \N__30999\
        );

    \I__5977\ : InMux
    port map (
            O => \N__31003\,
            I => \N__30996\
        );

    \I__5976\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30991\
        );

    \I__5975\ : Span4Mux_h
    port map (
            O => \N__30999\,
            I => \N__30986\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__30996\,
            I => \N__30986\
        );

    \I__5973\ : InMux
    port map (
            O => \N__30995\,
            I => \N__30983\
        );

    \I__5972\ : InMux
    port map (
            O => \N__30994\,
            I => \N__30980\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__30991\,
            I => \N__30975\
        );

    \I__5970\ : Span4Mux_v
    port map (
            O => \N__30986\,
            I => \N__30975\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__30983\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__30980\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5967\ : Odrv4
    port map (
            O => \N__30975\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5966\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30963\
        );

    \I__5965\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30960\
        );

    \I__5964\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30957\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__30963\,
            I => \N__30954\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__30960\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__30957\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__5960\ : Odrv12
    port map (
            O => \N__30954\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__5959\ : CascadeMux
    port map (
            O => \N__30947\,
            I => \N__30944\
        );

    \I__5958\ : InMux
    port map (
            O => \N__30944\,
            I => \N__30941\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__30941\,
            I => \N__30938\
        );

    \I__5956\ : Span4Mux_h
    port map (
            O => \N__30938\,
            I => \N__30935\
        );

    \I__5955\ : Span4Mux_v
    port map (
            O => \N__30935\,
            I => \N__30932\
        );

    \I__5954\ : Odrv4
    port map (
            O => \N__30932\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\
        );

    \I__5953\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30924\
        );

    \I__5952\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30921\
        );

    \I__5951\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30918\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__30924\,
            I => \N__30915\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__30921\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__30918\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__30915\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__5946\ : InMux
    port map (
            O => \N__30908\,
            I => \N__30904\
        );

    \I__5945\ : InMux
    port map (
            O => \N__30907\,
            I => \N__30901\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__30904\,
            I => \N__30897\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__30901\,
            I => \N__30894\
        );

    \I__5942\ : InMux
    port map (
            O => \N__30900\,
            I => \N__30889\
        );

    \I__5941\ : Span4Mux_v
    port map (
            O => \N__30897\,
            I => \N__30886\
        );

    \I__5940\ : Span12Mux_h
    port map (
            O => \N__30894\,
            I => \N__30883\
        );

    \I__5939\ : InMux
    port map (
            O => \N__30893\,
            I => \N__30880\
        );

    \I__5938\ : InMux
    port map (
            O => \N__30892\,
            I => \N__30877\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__30889\,
            I => \N__30872\
        );

    \I__5936\ : Span4Mux_v
    port map (
            O => \N__30886\,
            I => \N__30872\
        );

    \I__5935\ : Odrv12
    port map (
            O => \N__30883\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__30880\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__30877\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__30872\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5931\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30860\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__30860\,
            I => \N__30857\
        );

    \I__5929\ : Span4Mux_h
    port map (
            O => \N__30857\,
            I => \N__30854\
        );

    \I__5928\ : Odrv4
    port map (
            O => \N__30854\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__30851\,
            I => \N__30848\
        );

    \I__5926\ : InMux
    port map (
            O => \N__30848\,
            I => \N__30844\
        );

    \I__5925\ : InMux
    port map (
            O => \N__30847\,
            I => \N__30841\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__30844\,
            I => \N__30837\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__30841\,
            I => \N__30834\
        );

    \I__5922\ : InMux
    port map (
            O => \N__30840\,
            I => \N__30831\
        );

    \I__5921\ : Span4Mux_v
    port map (
            O => \N__30837\,
            I => \N__30826\
        );

    \I__5920\ : Span4Mux_v
    port map (
            O => \N__30834\,
            I => \N__30826\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__30831\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__30826\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__5917\ : InMux
    port map (
            O => \N__30821\,
            I => \N__30818\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__30818\,
            I => \N__30815\
        );

    \I__5915\ : Span4Mux_h
    port map (
            O => \N__30815\,
            I => \N__30812\
        );

    \I__5914\ : Odrv4
    port map (
            O => \N__30812\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\
        );

    \I__5913\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30805\
        );

    \I__5912\ : InMux
    port map (
            O => \N__30808\,
            I => \N__30801\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__30805\,
            I => \N__30798\
        );

    \I__5910\ : InMux
    port map (
            O => \N__30804\,
            I => \N__30795\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__30801\,
            I => \N__30792\
        );

    \I__5908\ : Span12Mux_h
    port map (
            O => \N__30798\,
            I => \N__30787\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__30795\,
            I => \N__30782\
        );

    \I__5906\ : Span4Mux_h
    port map (
            O => \N__30792\,
            I => \N__30782\
        );

    \I__5905\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30777\
        );

    \I__5904\ : InMux
    port map (
            O => \N__30790\,
            I => \N__30777\
        );

    \I__5903\ : Odrv12
    port map (
            O => \N__30787\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__5902\ : Odrv4
    port map (
            O => \N__30782\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__30777\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__5900\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30765\
        );

    \I__5899\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30762\
        );

    \I__5898\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30759\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__30765\,
            I => \N__30756\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__30762\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__30759\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5894\ : Odrv4
    port map (
            O => \N__30756\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5893\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30746\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__30746\,
            I => \N__30743\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__30743\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\
        );

    \I__5890\ : InMux
    port map (
            O => \N__30740\,
            I => \N__30735\
        );

    \I__5889\ : InMux
    port map (
            O => \N__30739\,
            I => \N__30732\
        );

    \I__5888\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30729\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__30735\,
            I => \N__30726\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__30732\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__30729\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__5884\ : Odrv12
    port map (
            O => \N__30726\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__5883\ : InMux
    port map (
            O => \N__30719\,
            I => \N__30716\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__30716\,
            I => \N__30713\
        );

    \I__5881\ : Span4Mux_h
    port map (
            O => \N__30713\,
            I => \N__30710\
        );

    \I__5880\ : Odrv4
    port map (
            O => \N__30710\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\
        );

    \I__5879\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30704\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__30704\,
            I => \N__30699\
        );

    \I__5877\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30696\
        );

    \I__5876\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30693\
        );

    \I__5875\ : Span4Mux_v
    port map (
            O => \N__30699\,
            I => \N__30690\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__30696\,
            I => \N__30687\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__30693\,
            I => \N__30682\
        );

    \I__5872\ : Span4Mux_h
    port map (
            O => \N__30690\,
            I => \N__30679\
        );

    \I__5871\ : Span4Mux_h
    port map (
            O => \N__30687\,
            I => \N__30676\
        );

    \I__5870\ : InMux
    port map (
            O => \N__30686\,
            I => \N__30671\
        );

    \I__5869\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30671\
        );

    \I__5868\ : Odrv4
    port map (
            O => \N__30682\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5867\ : Odrv4
    port map (
            O => \N__30679\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5866\ : Odrv4
    port map (
            O => \N__30676\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__30671\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5864\ : CascadeMux
    port map (
            O => \N__30662\,
            I => \N__30659\
        );

    \I__5863\ : InMux
    port map (
            O => \N__30659\,
            I => \N__30656\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__30656\,
            I => \N__30653\
        );

    \I__5861\ : Span4Mux_h
    port map (
            O => \N__30653\,
            I => \N__30650\
        );

    \I__5860\ : Odrv4
    port map (
            O => \N__30650\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\
        );

    \I__5859\ : CascadeMux
    port map (
            O => \N__30647\,
            I => \N__30644\
        );

    \I__5858\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30640\
        );

    \I__5857\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30637\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__30640\,
            I => \N__30634\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__30637\,
            I => \N__30631\
        );

    \I__5854\ : Span4Mux_v
    port map (
            O => \N__30634\,
            I => \N__30627\
        );

    \I__5853\ : Span4Mux_h
    port map (
            O => \N__30631\,
            I => \N__30622\
        );

    \I__5852\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30619\
        );

    \I__5851\ : Span4Mux_h
    port map (
            O => \N__30627\,
            I => \N__30616\
        );

    \I__5850\ : InMux
    port map (
            O => \N__30626\,
            I => \N__30611\
        );

    \I__5849\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30611\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__30622\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__30619\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__5846\ : Odrv4
    port map (
            O => \N__30616\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__30611\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__5844\ : InMux
    port map (
            O => \N__30602\,
            I => \N__30599\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__30599\,
            I => \N__30596\
        );

    \I__5842\ : Span4Mux_h
    port map (
            O => \N__30596\,
            I => \N__30591\
        );

    \I__5841\ : CascadeMux
    port map (
            O => \N__30595\,
            I => \N__30588\
        );

    \I__5840\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30585\
        );

    \I__5839\ : Span4Mux_v
    port map (
            O => \N__30591\,
            I => \N__30582\
        );

    \I__5838\ : InMux
    port map (
            O => \N__30588\,
            I => \N__30579\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__30585\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__5836\ : Odrv4
    port map (
            O => \N__30582\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__30579\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__5834\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30569\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__30569\,
            I => \N__30566\
        );

    \I__5832\ : Span4Mux_v
    port map (
            O => \N__30566\,
            I => \N__30563\
        );

    \I__5831\ : Odrv4
    port map (
            O => \N__30563\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\
        );

    \I__5830\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30555\
        );

    \I__5829\ : InMux
    port map (
            O => \N__30559\,
            I => \N__30552\
        );

    \I__5828\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30549\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__30555\,
            I => \N__30546\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__30552\,
            I => \N__30543\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__30549\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5824\ : Odrv4
    port map (
            O => \N__30546\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5823\ : Odrv12
    port map (
            O => \N__30543\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__30536\,
            I => \N__30533\
        );

    \I__5821\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30530\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__30530\,
            I => \N__30525\
        );

    \I__5819\ : InMux
    port map (
            O => \N__30529\,
            I => \N__30520\
        );

    \I__5818\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30517\
        );

    \I__5817\ : Span4Mux_v
    port map (
            O => \N__30525\,
            I => \N__30514\
        );

    \I__5816\ : CascadeMux
    port map (
            O => \N__30524\,
            I => \N__30511\
        );

    \I__5815\ : CascadeMux
    port map (
            O => \N__30523\,
            I => \N__30508\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__30520\,
            I => \N__30505\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__30517\,
            I => \N__30502\
        );

    \I__5812\ : Span4Mux_h
    port map (
            O => \N__30514\,
            I => \N__30499\
        );

    \I__5811\ : InMux
    port map (
            O => \N__30511\,
            I => \N__30496\
        );

    \I__5810\ : InMux
    port map (
            O => \N__30508\,
            I => \N__30493\
        );

    \I__5809\ : Span4Mux_h
    port map (
            O => \N__30505\,
            I => \N__30490\
        );

    \I__5808\ : Odrv12
    port map (
            O => \N__30502\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5807\ : Odrv4
    port map (
            O => \N__30499\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__30496\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__30493\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5804\ : Odrv4
    port map (
            O => \N__30490\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5803\ : CascadeMux
    port map (
            O => \N__30479\,
            I => \N__30476\
        );

    \I__5802\ : InMux
    port map (
            O => \N__30476\,
            I => \N__30473\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__30473\,
            I => \N__30470\
        );

    \I__5800\ : Span4Mux_h
    port map (
            O => \N__30470\,
            I => \N__30467\
        );

    \I__5799\ : Odrv4
    port map (
            O => \N__30467\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\
        );

    \I__5798\ : InMux
    port map (
            O => \N__30464\,
            I => \N__30459\
        );

    \I__5797\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30456\
        );

    \I__5796\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30453\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__30459\,
            I => \N__30450\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__30456\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__30453\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__5792\ : Odrv12
    port map (
            O => \N__30450\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__5791\ : CascadeMux
    port map (
            O => \N__30443\,
            I => \N__30440\
        );

    \I__5790\ : InMux
    port map (
            O => \N__30440\,
            I => \N__30436\
        );

    \I__5789\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30433\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__30436\,
            I => \N__30429\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__30433\,
            I => \N__30426\
        );

    \I__5786\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30423\
        );

    \I__5785\ : Span4Mux_v
    port map (
            O => \N__30429\,
            I => \N__30418\
        );

    \I__5784\ : Span4Mux_h
    port map (
            O => \N__30426\,
            I => \N__30413\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__30423\,
            I => \N__30413\
        );

    \I__5782\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30410\
        );

    \I__5781\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30407\
        );

    \I__5780\ : Span4Mux_h
    port map (
            O => \N__30418\,
            I => \N__30404\
        );

    \I__5779\ : Span4Mux_h
    port map (
            O => \N__30413\,
            I => \N__30399\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__30410\,
            I => \N__30399\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__30407\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__5776\ : Odrv4
    port map (
            O => \N__30404\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__5775\ : Odrv4
    port map (
            O => \N__30399\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__5774\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30389\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__30389\,
            I => \N__30386\
        );

    \I__5772\ : Odrv4
    port map (
            O => \N__30386\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\
        );

    \I__5771\ : InMux
    port map (
            O => \N__30383\,
            I => \N__30379\
        );

    \I__5770\ : InMux
    port map (
            O => \N__30382\,
            I => \N__30376\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__30379\,
            I => \N__30373\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__30376\,
            I => \N__30370\
        );

    \I__5767\ : Span12Mux_h
    port map (
            O => \N__30373\,
            I => \N__30364\
        );

    \I__5766\ : Span4Mux_h
    port map (
            O => \N__30370\,
            I => \N__30361\
        );

    \I__5765\ : InMux
    port map (
            O => \N__30369\,
            I => \N__30358\
        );

    \I__5764\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30353\
        );

    \I__5763\ : InMux
    port map (
            O => \N__30367\,
            I => \N__30353\
        );

    \I__5762\ : Odrv12
    port map (
            O => \N__30364\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__30361\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__30358\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__30353\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__30344\,
            I => \N__30341\
        );

    \I__5757\ : InMux
    port map (
            O => \N__30341\,
            I => \N__30338\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__30338\,
            I => \N__30335\
        );

    \I__5755\ : Span4Mux_v
    port map (
            O => \N__30335\,
            I => \N__30331\
        );

    \I__5754\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30327\
        );

    \I__5753\ : Span4Mux_v
    port map (
            O => \N__30331\,
            I => \N__30324\
        );

    \I__5752\ : InMux
    port map (
            O => \N__30330\,
            I => \N__30321\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__30327\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__30324\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__30321\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5748\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30311\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__30311\,
            I => \N__30308\
        );

    \I__5746\ : Span4Mux_v
    port map (
            O => \N__30308\,
            I => \N__30305\
        );

    \I__5745\ : Odrv4
    port map (
            O => \N__30305\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_8\
        );

    \I__5744\ : InMux
    port map (
            O => \N__30302\,
            I => \N__30298\
        );

    \I__5743\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30295\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__30298\,
            I => \N__30291\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__30295\,
            I => \N__30288\
        );

    \I__5740\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30283\
        );

    \I__5739\ : Span12Mux_v
    port map (
            O => \N__30291\,
            I => \N__30280\
        );

    \I__5738\ : Span4Mux_v
    port map (
            O => \N__30288\,
            I => \N__30277\
        );

    \I__5737\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30272\
        );

    \I__5736\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30272\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__30283\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__5734\ : Odrv12
    port map (
            O => \N__30280\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__5733\ : Odrv4
    port map (
            O => \N__30277\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__30272\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__5731\ : InMux
    port map (
            O => \N__30263\,
            I => \N__30260\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__30260\,
            I => \N__30257\
        );

    \I__5729\ : Span4Mux_h
    port map (
            O => \N__30257\,
            I => \N__30254\
        );

    \I__5728\ : Odrv4
    port map (
            O => \N__30254\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30246\
        );

    \I__5726\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30243\
        );

    \I__5725\ : InMux
    port map (
            O => \N__30249\,
            I => \N__30240\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__30246\,
            I => \N__30237\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__30243\,
            I => \N__30234\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__30240\,
            I => \N__30231\
        );

    \I__5721\ : Span4Mux_h
    port map (
            O => \N__30237\,
            I => \N__30228\
        );

    \I__5720\ : Span4Mux_v
    port map (
            O => \N__30234\,
            I => \N__30223\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__30231\,
            I => \N__30223\
        );

    \I__5718\ : Odrv4
    port map (
            O => \N__30228\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__30223\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5716\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30215\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__30215\,
            I => \N__30212\
        );

    \I__5714\ : Span4Mux_h
    port map (
            O => \N__30212\,
            I => \N__30209\
        );

    \I__5713\ : Odrv4
    port map (
            O => \N__30209\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_11\
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__30206\,
            I => \N__30203\
        );

    \I__5711\ : InMux
    port map (
            O => \N__30203\,
            I => \N__30198\
        );

    \I__5710\ : InMux
    port map (
            O => \N__30202\,
            I => \N__30195\
        );

    \I__5709\ : InMux
    port map (
            O => \N__30201\,
            I => \N__30192\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__30198\,
            I => \N__30187\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__30195\,
            I => \N__30187\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__30192\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__5705\ : Odrv12
    port map (
            O => \N__30187\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__5704\ : InMux
    port map (
            O => \N__30182\,
            I => \bfn_13_27_0_\
        );

    \I__5703\ : CascadeMux
    port map (
            O => \N__30179\,
            I => \N__30176\
        );

    \I__5702\ : InMux
    port map (
            O => \N__30176\,
            I => \N__30172\
        );

    \I__5701\ : InMux
    port map (
            O => \N__30175\,
            I => \N__30169\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__30172\,
            I => \N__30163\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__30169\,
            I => \N__30163\
        );

    \I__5698\ : InMux
    port map (
            O => \N__30168\,
            I => \N__30160\
        );

    \I__5697\ : Span4Mux_v
    port map (
            O => \N__30163\,
            I => \N__30157\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__30160\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__5695\ : Odrv4
    port map (
            O => \N__30157\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__5694\ : InMux
    port map (
            O => \N__30152\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__5693\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30143\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30143\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__30143\,
            I => \N__30139\
        );

    \I__5690\ : InMux
    port map (
            O => \N__30142\,
            I => \N__30136\
        );

    \I__5689\ : Span4Mux_v
    port map (
            O => \N__30139\,
            I => \N__30133\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__30136\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__5687\ : Odrv4
    port map (
            O => \N__30133\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__5686\ : InMux
    port map (
            O => \N__30128\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__5685\ : InMux
    port map (
            O => \N__30125\,
            I => \N__30118\
        );

    \I__5684\ : InMux
    port map (
            O => \N__30124\,
            I => \N__30118\
        );

    \I__5683\ : InMux
    port map (
            O => \N__30123\,
            I => \N__30115\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__30118\,
            I => \N__30112\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__30115\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__5680\ : Odrv12
    port map (
            O => \N__30112\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__5679\ : InMux
    port map (
            O => \N__30107\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__30104\,
            I => \N__30101\
        );

    \I__5677\ : InMux
    port map (
            O => \N__30101\,
            I => \N__30098\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__30098\,
            I => \N__30094\
        );

    \I__5675\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30091\
        );

    \I__5674\ : Span4Mux_v
    port map (
            O => \N__30094\,
            I => \N__30088\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__30091\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__30088\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__5671\ : InMux
    port map (
            O => \N__30083\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__5670\ : InMux
    port map (
            O => \N__30080\,
            I => \N__30060\
        );

    \I__5669\ : InMux
    port map (
            O => \N__30079\,
            I => \N__30060\
        );

    \I__5668\ : InMux
    port map (
            O => \N__30078\,
            I => \N__30060\
        );

    \I__5667\ : InMux
    port map (
            O => \N__30077\,
            I => \N__30060\
        );

    \I__5666\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30033\
        );

    \I__5665\ : InMux
    port map (
            O => \N__30075\,
            I => \N__30033\
        );

    \I__5664\ : InMux
    port map (
            O => \N__30074\,
            I => \N__30033\
        );

    \I__5663\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30033\
        );

    \I__5662\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30024\
        );

    \I__5661\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30024\
        );

    \I__5660\ : InMux
    port map (
            O => \N__30070\,
            I => \N__30024\
        );

    \I__5659\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30024\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__30060\,
            I => \N__30021\
        );

    \I__5657\ : InMux
    port map (
            O => \N__30059\,
            I => \N__30016\
        );

    \I__5656\ : InMux
    port map (
            O => \N__30058\,
            I => \N__30016\
        );

    \I__5655\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30007\
        );

    \I__5654\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30007\
        );

    \I__5653\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30007\
        );

    \I__5652\ : InMux
    port map (
            O => \N__30054\,
            I => \N__30007\
        );

    \I__5651\ : InMux
    port map (
            O => \N__30053\,
            I => \N__29998\
        );

    \I__5650\ : InMux
    port map (
            O => \N__30052\,
            I => \N__29998\
        );

    \I__5649\ : InMux
    port map (
            O => \N__30051\,
            I => \N__29998\
        );

    \I__5648\ : InMux
    port map (
            O => \N__30050\,
            I => \N__29998\
        );

    \I__5647\ : InMux
    port map (
            O => \N__30049\,
            I => \N__29989\
        );

    \I__5646\ : InMux
    port map (
            O => \N__30048\,
            I => \N__29989\
        );

    \I__5645\ : InMux
    port map (
            O => \N__30047\,
            I => \N__29989\
        );

    \I__5644\ : InMux
    port map (
            O => \N__30046\,
            I => \N__29989\
        );

    \I__5643\ : InMux
    port map (
            O => \N__30045\,
            I => \N__29980\
        );

    \I__5642\ : InMux
    port map (
            O => \N__30044\,
            I => \N__29980\
        );

    \I__5641\ : InMux
    port map (
            O => \N__30043\,
            I => \N__29980\
        );

    \I__5640\ : InMux
    port map (
            O => \N__30042\,
            I => \N__29980\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__30033\,
            I => \N__29975\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__30024\,
            I => \N__29975\
        );

    \I__5637\ : Odrv4
    port map (
            O => \N__30021\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__30016\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__30007\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__29998\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__29989\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__29980\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__5631\ : Odrv4
    port map (
            O => \N__29975\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__5630\ : InMux
    port map (
            O => \N__29960\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__5629\ : CascadeMux
    port map (
            O => \N__29957\,
            I => \N__29954\
        );

    \I__5628\ : InMux
    port map (
            O => \N__29954\,
            I => \N__29951\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__29951\,
            I => \N__29947\
        );

    \I__5626\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29944\
        );

    \I__5625\ : Span4Mux_v
    port map (
            O => \N__29947\,
            I => \N__29941\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__29944\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__5623\ : Odrv4
    port map (
            O => \N__29941\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__5622\ : CEMux
    port map (
            O => \N__29936\,
            I => \N__29933\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__29933\,
            I => \N__29927\
        );

    \I__5620\ : CEMux
    port map (
            O => \N__29932\,
            I => \N__29924\
        );

    \I__5619\ : CEMux
    port map (
            O => \N__29931\,
            I => \N__29921\
        );

    \I__5618\ : CEMux
    port map (
            O => \N__29930\,
            I => \N__29918\
        );

    \I__5617\ : Span4Mux_h
    port map (
            O => \N__29927\,
            I => \N__29915\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__29924\,
            I => \N__29910\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__29921\,
            I => \N__29910\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__29918\,
            I => \N__29907\
        );

    \I__5613\ : Odrv4
    port map (
            O => \N__29915\,
            I => \current_shift_inst.timer_s1.N_167_i\
        );

    \I__5612\ : Odrv4
    port map (
            O => \N__29910\,
            I => \current_shift_inst.timer_s1.N_167_i\
        );

    \I__5611\ : Odrv4
    port map (
            O => \N__29907\,
            I => \current_shift_inst.timer_s1.N_167_i\
        );

    \I__5610\ : InMux
    port map (
            O => \N__29900\,
            I => \N__29894\
        );

    \I__5609\ : InMux
    port map (
            O => \N__29899\,
            I => \N__29894\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__29894\,
            I => \N__29890\
        );

    \I__5607\ : InMux
    port map (
            O => \N__29893\,
            I => \N__29887\
        );

    \I__5606\ : Span4Mux_v
    port map (
            O => \N__29890\,
            I => \N__29884\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__29887\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__5604\ : Odrv4
    port map (
            O => \N__29884\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__5603\ : InMux
    port map (
            O => \N__29879\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__5602\ : CascadeMux
    port map (
            O => \N__29876\,
            I => \N__29873\
        );

    \I__5601\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29869\
        );

    \I__5600\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29866\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__29869\,
            I => \N__29862\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29859\
        );

    \I__5597\ : InMux
    port map (
            O => \N__29865\,
            I => \N__29856\
        );

    \I__5596\ : Span4Mux_v
    port map (
            O => \N__29862\,
            I => \N__29851\
        );

    \I__5595\ : Span4Mux_v
    port map (
            O => \N__29859\,
            I => \N__29851\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__29856\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__29851\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__5592\ : InMux
    port map (
            O => \N__29846\,
            I => \bfn_13_26_0_\
        );

    \I__5591\ : CascadeMux
    port map (
            O => \N__29843\,
            I => \N__29839\
        );

    \I__5590\ : CascadeMux
    port map (
            O => \N__29842\,
            I => \N__29836\
        );

    \I__5589\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29833\
        );

    \I__5588\ : InMux
    port map (
            O => \N__29836\,
            I => \N__29830\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__29833\,
            I => \N__29826\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__29830\,
            I => \N__29823\
        );

    \I__5585\ : InMux
    port map (
            O => \N__29829\,
            I => \N__29820\
        );

    \I__5584\ : Span4Mux_v
    port map (
            O => \N__29826\,
            I => \N__29815\
        );

    \I__5583\ : Span4Mux_v
    port map (
            O => \N__29823\,
            I => \N__29815\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__29820\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__5581\ : Odrv4
    port map (
            O => \N__29815\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__5580\ : InMux
    port map (
            O => \N__29810\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__5579\ : InMux
    port map (
            O => \N__29807\,
            I => \N__29801\
        );

    \I__5578\ : InMux
    port map (
            O => \N__29806\,
            I => \N__29801\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__29801\,
            I => \N__29797\
        );

    \I__5576\ : InMux
    port map (
            O => \N__29800\,
            I => \N__29794\
        );

    \I__5575\ : Span4Mux_v
    port map (
            O => \N__29797\,
            I => \N__29791\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__29794\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__29791\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__5572\ : InMux
    port map (
            O => \N__29786\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__5571\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29776\
        );

    \I__5570\ : InMux
    port map (
            O => \N__29782\,
            I => \N__29776\
        );

    \I__5569\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29773\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__29776\,
            I => \N__29770\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__29773\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__5566\ : Odrv12
    port map (
            O => \N__29770\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__5565\ : InMux
    port map (
            O => \N__29765\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__5564\ : CascadeMux
    port map (
            O => \N__29762\,
            I => \N__29758\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__29761\,
            I => \N__29755\
        );

    \I__5562\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29750\
        );

    \I__5561\ : InMux
    port map (
            O => \N__29755\,
            I => \N__29750\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__29750\,
            I => \N__29746\
        );

    \I__5559\ : InMux
    port map (
            O => \N__29749\,
            I => \N__29743\
        );

    \I__5558\ : Span4Mux_v
    port map (
            O => \N__29746\,
            I => \N__29740\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__29743\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__5556\ : Odrv4
    port map (
            O => \N__29740\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__5555\ : InMux
    port map (
            O => \N__29735\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__5554\ : CascadeMux
    port map (
            O => \N__29732\,
            I => \N__29728\
        );

    \I__5553\ : CascadeMux
    port map (
            O => \N__29731\,
            I => \N__29725\
        );

    \I__5552\ : InMux
    port map (
            O => \N__29728\,
            I => \N__29720\
        );

    \I__5551\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29720\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__29720\,
            I => \N__29716\
        );

    \I__5549\ : InMux
    port map (
            O => \N__29719\,
            I => \N__29713\
        );

    \I__5548\ : Span4Mux_v
    port map (
            O => \N__29716\,
            I => \N__29710\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__29713\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__5546\ : Odrv4
    port map (
            O => \N__29710\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__5545\ : InMux
    port map (
            O => \N__29705\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__29702\,
            I => \N__29699\
        );

    \I__5543\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29694\
        );

    \I__5542\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29691\
        );

    \I__5541\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29688\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__29694\,
            I => \N__29683\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__29691\,
            I => \N__29683\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__29688\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__5537\ : Odrv12
    port map (
            O => \N__29683\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__5536\ : InMux
    port map (
            O => \N__29678\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__5535\ : CascadeMux
    port map (
            O => \N__29675\,
            I => \N__29672\
        );

    \I__5534\ : InMux
    port map (
            O => \N__29672\,
            I => \N__29668\
        );

    \I__5533\ : InMux
    port map (
            O => \N__29671\,
            I => \N__29665\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__29668\,
            I => \N__29659\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__29665\,
            I => \N__29659\
        );

    \I__5530\ : InMux
    port map (
            O => \N__29664\,
            I => \N__29656\
        );

    \I__5529\ : Span4Mux_v
    port map (
            O => \N__29659\,
            I => \N__29653\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__29656\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__5527\ : Odrv4
    port map (
            O => \N__29653\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__5526\ : InMux
    port map (
            O => \N__29648\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__5525\ : InMux
    port map (
            O => \N__29645\,
            I => \N__29639\
        );

    \I__5524\ : InMux
    port map (
            O => \N__29644\,
            I => \N__29639\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__29639\,
            I => \N__29635\
        );

    \I__5522\ : InMux
    port map (
            O => \N__29638\,
            I => \N__29632\
        );

    \I__5521\ : Span4Mux_v
    port map (
            O => \N__29635\,
            I => \N__29629\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__29632\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__5519\ : Odrv4
    port map (
            O => \N__29629\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__5518\ : InMux
    port map (
            O => \N__29624\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__5517\ : CascadeMux
    port map (
            O => \N__29621\,
            I => \N__29618\
        );

    \I__5516\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29615\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__29615\,
            I => \N__29610\
        );

    \I__5514\ : InMux
    port map (
            O => \N__29614\,
            I => \N__29607\
        );

    \I__5513\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29604\
        );

    \I__5512\ : Span4Mux_v
    port map (
            O => \N__29610\,
            I => \N__29601\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__29607\,
            I => \N__29598\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__29604\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__5509\ : Odrv4
    port map (
            O => \N__29601\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__5508\ : Odrv12
    port map (
            O => \N__29598\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__5507\ : InMux
    port map (
            O => \N__29591\,
            I => \bfn_13_25_0_\
        );

    \I__5506\ : CascadeMux
    port map (
            O => \N__29588\,
            I => \N__29585\
        );

    \I__5505\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29581\
        );

    \I__5504\ : CascadeMux
    port map (
            O => \N__29584\,
            I => \N__29578\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__29581\,
            I => \N__29574\
        );

    \I__5502\ : InMux
    port map (
            O => \N__29578\,
            I => \N__29571\
        );

    \I__5501\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29568\
        );

    \I__5500\ : Span4Mux_v
    port map (
            O => \N__29574\,
            I => \N__29565\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__29571\,
            I => \N__29562\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__29568\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__29565\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__5496\ : Odrv12
    port map (
            O => \N__29562\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__5495\ : InMux
    port map (
            O => \N__29555\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__5494\ : InMux
    port map (
            O => \N__29552\,
            I => \N__29546\
        );

    \I__5493\ : InMux
    port map (
            O => \N__29551\,
            I => \N__29546\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__29546\,
            I => \N__29542\
        );

    \I__5491\ : InMux
    port map (
            O => \N__29545\,
            I => \N__29539\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__29542\,
            I => \N__29536\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__29539\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__29536\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__5487\ : InMux
    port map (
            O => \N__29531\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__5486\ : InMux
    port map (
            O => \N__29528\,
            I => \N__29521\
        );

    \I__5485\ : InMux
    port map (
            O => \N__29527\,
            I => \N__29521\
        );

    \I__5484\ : InMux
    port map (
            O => \N__29526\,
            I => \N__29518\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__29521\,
            I => \N__29515\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__29518\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__5481\ : Odrv12
    port map (
            O => \N__29515\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__5480\ : InMux
    port map (
            O => \N__29510\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__5479\ : CascadeMux
    port map (
            O => \N__29507\,
            I => \N__29503\
        );

    \I__5478\ : CascadeMux
    port map (
            O => \N__29506\,
            I => \N__29500\
        );

    \I__5477\ : InMux
    port map (
            O => \N__29503\,
            I => \N__29495\
        );

    \I__5476\ : InMux
    port map (
            O => \N__29500\,
            I => \N__29495\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__29495\,
            I => \N__29491\
        );

    \I__5474\ : InMux
    port map (
            O => \N__29494\,
            I => \N__29488\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__29491\,
            I => \N__29485\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__29488\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__29485\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__5470\ : InMux
    port map (
            O => \N__29480\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__5469\ : CascadeMux
    port map (
            O => \N__29477\,
            I => \N__29473\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__29476\,
            I => \N__29470\
        );

    \I__5467\ : InMux
    port map (
            O => \N__29473\,
            I => \N__29465\
        );

    \I__5466\ : InMux
    port map (
            O => \N__29470\,
            I => \N__29465\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__29465\,
            I => \N__29461\
        );

    \I__5464\ : InMux
    port map (
            O => \N__29464\,
            I => \N__29458\
        );

    \I__5463\ : Span4Mux_v
    port map (
            O => \N__29461\,
            I => \N__29455\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__29458\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__29455\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__5460\ : InMux
    port map (
            O => \N__29450\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__5459\ : CascadeMux
    port map (
            O => \N__29447\,
            I => \N__29444\
        );

    \I__5458\ : InMux
    port map (
            O => \N__29444\,
            I => \N__29440\
        );

    \I__5457\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29437\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__29440\,
            I => \N__29431\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__29437\,
            I => \N__29431\
        );

    \I__5454\ : InMux
    port map (
            O => \N__29436\,
            I => \N__29428\
        );

    \I__5453\ : Span4Mux_v
    port map (
            O => \N__29431\,
            I => \N__29425\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__29428\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__5451\ : Odrv4
    port map (
            O => \N__29425\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__5450\ : InMux
    port map (
            O => \N__29420\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__5449\ : InMux
    port map (
            O => \N__29417\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__5448\ : InMux
    port map (
            O => \N__29414\,
            I => \N__29407\
        );

    \I__5447\ : InMux
    port map (
            O => \N__29413\,
            I => \N__29407\
        );

    \I__5446\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29404\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__29407\,
            I => \N__29400\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__29404\,
            I => \N__29397\
        );

    \I__5443\ : InMux
    port map (
            O => \N__29403\,
            I => \N__29394\
        );

    \I__5442\ : Span4Mux_v
    port map (
            O => \N__29400\,
            I => \N__29391\
        );

    \I__5441\ : Odrv12
    port map (
            O => \N__29397\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__29394\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__29391\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__5438\ : IoInMux
    port map (
            O => \N__29384\,
            I => \N__29381\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__29381\,
            I => \N__29378\
        );

    \I__5436\ : Odrv12
    port map (
            O => \N__29378\,
            I => s2_phy_c
        );

    \I__5435\ : InMux
    port map (
            O => \N__29375\,
            I => \bfn_13_24_0_\
        );

    \I__5434\ : InMux
    port map (
            O => \N__29372\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__5433\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29362\
        );

    \I__5432\ : InMux
    port map (
            O => \N__29368\,
            I => \N__29362\
        );

    \I__5431\ : InMux
    port map (
            O => \N__29367\,
            I => \N__29359\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__29362\,
            I => \N__29356\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__29359\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__5428\ : Odrv12
    port map (
            O => \N__29356\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__5427\ : InMux
    port map (
            O => \N__29351\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__5426\ : CascadeMux
    port map (
            O => \N__29348\,
            I => \N__29344\
        );

    \I__5425\ : InMux
    port map (
            O => \N__29347\,
            I => \N__29340\
        );

    \I__5424\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29337\
        );

    \I__5423\ : InMux
    port map (
            O => \N__29343\,
            I => \N__29334\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__29340\,
            I => \N__29327\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__29337\,
            I => \N__29327\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__29334\,
            I => \N__29327\
        );

    \I__5419\ : Odrv12
    port map (
            O => \N__29327\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__5418\ : InMux
    port map (
            O => \N__29324\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__5417\ : CascadeMux
    port map (
            O => \N__29321\,
            I => \N__29317\
        );

    \I__5416\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29314\
        );

    \I__5415\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29311\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__29314\,
            I => \N__29305\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__29311\,
            I => \N__29305\
        );

    \I__5412\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29302\
        );

    \I__5411\ : Span4Mux_v
    port map (
            O => \N__29305\,
            I => \N__29299\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__29302\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__5409\ : Odrv4
    port map (
            O => \N__29299\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__5408\ : InMux
    port map (
            O => \N__29294\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__29291\,
            I => \N__29288\
        );

    \I__5406\ : InMux
    port map (
            O => \N__29288\,
            I => \N__29284\
        );

    \I__5405\ : InMux
    port map (
            O => \N__29287\,
            I => \N__29281\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__29284\,
            I => \N__29275\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__29281\,
            I => \N__29275\
        );

    \I__5402\ : InMux
    port map (
            O => \N__29280\,
            I => \N__29272\
        );

    \I__5401\ : Span4Mux_v
    port map (
            O => \N__29275\,
            I => \N__29269\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__29272\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__5399\ : Odrv4
    port map (
            O => \N__29269\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__5398\ : InMux
    port map (
            O => \N__29264\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__29261\,
            I => \N__29257\
        );

    \I__5396\ : CascadeMux
    port map (
            O => \N__29260\,
            I => \N__29254\
        );

    \I__5395\ : InMux
    port map (
            O => \N__29257\,
            I => \N__29249\
        );

    \I__5394\ : InMux
    port map (
            O => \N__29254\,
            I => \N__29249\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__29249\,
            I => \N__29245\
        );

    \I__5392\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29242\
        );

    \I__5391\ : Span4Mux_v
    port map (
            O => \N__29245\,
            I => \N__29239\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__29242\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__5389\ : Odrv4
    port map (
            O => \N__29239\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__5388\ : InMux
    port map (
            O => \N__29234\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__5387\ : InMux
    port map (
            O => \N__29231\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__5386\ : InMux
    port map (
            O => \N__29228\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__5385\ : InMux
    port map (
            O => \N__29225\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__5384\ : InMux
    port map (
            O => \N__29222\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__5383\ : InMux
    port map (
            O => \N__29219\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__5382\ : InMux
    port map (
            O => \N__29216\,
            I => \bfn_13_22_0_\
        );

    \I__5381\ : InMux
    port map (
            O => \N__29213\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__5380\ : InMux
    port map (
            O => \N__29210\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__5379\ : InMux
    port map (
            O => \N__29207\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__5378\ : InMux
    port map (
            O => \N__29204\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__5377\ : InMux
    port map (
            O => \N__29201\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__5376\ : InMux
    port map (
            O => \N__29198\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__5375\ : InMux
    port map (
            O => \N__29195\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__5374\ : InMux
    port map (
            O => \N__29192\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__5373\ : InMux
    port map (
            O => \N__29189\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__5372\ : InMux
    port map (
            O => \N__29186\,
            I => \bfn_13_21_0_\
        );

    \I__5371\ : InMux
    port map (
            O => \N__29183\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__5370\ : InMux
    port map (
            O => \N__29180\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__5369\ : InMux
    port map (
            O => \N__29177\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__5368\ : InMux
    port map (
            O => \N__29174\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__5367\ : InMux
    port map (
            O => \N__29171\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__5366\ : InMux
    port map (
            O => \N__29168\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__5365\ : InMux
    port map (
            O => \N__29165\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__5364\ : InMux
    port map (
            O => \N__29162\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__5363\ : InMux
    port map (
            O => \N__29159\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__5362\ : InMux
    port map (
            O => \N__29156\,
            I => \bfn_13_20_0_\
        );

    \I__5361\ : InMux
    port map (
            O => \N__29153\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__5360\ : InMux
    port map (
            O => \N__29150\,
            I => \N__29147\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__29147\,
            I => \current_shift_inst.un38_control_input_cry_1_c_RNOZ0\
        );

    \I__5358\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29140\
        );

    \I__5357\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29137\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__29140\,
            I => \N__29132\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__29137\,
            I => \N__29129\
        );

    \I__5354\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29126\
        );

    \I__5353\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29123\
        );

    \I__5352\ : Span12Mux_v
    port map (
            O => \N__29132\,
            I => \N__29120\
        );

    \I__5351\ : Span12Mux_v
    port map (
            O => \N__29129\,
            I => \N__29117\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__29126\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__29123\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5348\ : Odrv12
    port map (
            O => \N__29120\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5347\ : Odrv12
    port map (
            O => \N__29117\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5346\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29105\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__29105\,
            I => \N__29101\
        );

    \I__5344\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29098\
        );

    \I__5343\ : Span4Mux_v
    port map (
            O => \N__29101\,
            I => \N__29094\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29091\
        );

    \I__5341\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29088\
        );

    \I__5340\ : Span4Mux_h
    port map (
            O => \N__29094\,
            I => \N__29083\
        );

    \I__5339\ : Span4Mux_v
    port map (
            O => \N__29091\,
            I => \N__29083\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__29088\,
            I => \N__29080\
        );

    \I__5337\ : Span4Mux_v
    port map (
            O => \N__29083\,
            I => \N__29077\
        );

    \I__5336\ : Span12Mux_v
    port map (
            O => \N__29080\,
            I => \N__29074\
        );

    \I__5335\ : Span4Mux_v
    port map (
            O => \N__29077\,
            I => \N__29071\
        );

    \I__5334\ : Odrv12
    port map (
            O => \N__29074\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__29071\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__5332\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29062\
        );

    \I__5331\ : InMux
    port map (
            O => \N__29065\,
            I => \N__29059\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__29062\,
            I => \N__29056\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__29059\,
            I => \N__29051\
        );

    \I__5328\ : Span4Mux_v
    port map (
            O => \N__29056\,
            I => \N__29048\
        );

    \I__5327\ : InMux
    port map (
            O => \N__29055\,
            I => \N__29043\
        );

    \I__5326\ : InMux
    port map (
            O => \N__29054\,
            I => \N__29043\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__29051\,
            I => \N__29040\
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__29048\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__29043\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__29040\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5321\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29021\
        );

    \I__5320\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29021\
        );

    \I__5319\ : InMux
    port map (
            O => \N__29031\,
            I => \N__29021\
        );

    \I__5318\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29021\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__29021\,
            I => \N__28996\
        );

    \I__5316\ : InMux
    port map (
            O => \N__29020\,
            I => \N__28987\
        );

    \I__5315\ : InMux
    port map (
            O => \N__29019\,
            I => \N__28987\
        );

    \I__5314\ : InMux
    port map (
            O => \N__29018\,
            I => \N__28987\
        );

    \I__5313\ : InMux
    port map (
            O => \N__29017\,
            I => \N__28987\
        );

    \I__5312\ : InMux
    port map (
            O => \N__29016\,
            I => \N__28978\
        );

    \I__5311\ : InMux
    port map (
            O => \N__29015\,
            I => \N__28978\
        );

    \I__5310\ : InMux
    port map (
            O => \N__29014\,
            I => \N__28978\
        );

    \I__5309\ : InMux
    port map (
            O => \N__29013\,
            I => \N__28978\
        );

    \I__5308\ : InMux
    port map (
            O => \N__29012\,
            I => \N__28969\
        );

    \I__5307\ : InMux
    port map (
            O => \N__29011\,
            I => \N__28969\
        );

    \I__5306\ : InMux
    port map (
            O => \N__29010\,
            I => \N__28960\
        );

    \I__5305\ : InMux
    port map (
            O => \N__29009\,
            I => \N__28960\
        );

    \I__5304\ : InMux
    port map (
            O => \N__29008\,
            I => \N__28960\
        );

    \I__5303\ : InMux
    port map (
            O => \N__29007\,
            I => \N__28960\
        );

    \I__5302\ : InMux
    port map (
            O => \N__29006\,
            I => \N__28951\
        );

    \I__5301\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28951\
        );

    \I__5300\ : InMux
    port map (
            O => \N__29004\,
            I => \N__28951\
        );

    \I__5299\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28951\
        );

    \I__5298\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28942\
        );

    \I__5297\ : InMux
    port map (
            O => \N__29001\,
            I => \N__28942\
        );

    \I__5296\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28942\
        );

    \I__5295\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28942\
        );

    \I__5294\ : Span4Mux_v
    port map (
            O => \N__28996\,
            I => \N__28935\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__28987\,
            I => \N__28935\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__28978\,
            I => \N__28935\
        );

    \I__5291\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28926\
        );

    \I__5290\ : InMux
    port map (
            O => \N__28976\,
            I => \N__28926\
        );

    \I__5289\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28926\
        );

    \I__5288\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28926\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__28969\,
            I => \N__28921\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__28960\,
            I => \N__28921\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28918\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__28942\,
            I => \N__28913\
        );

    \I__5283\ : Span4Mux_v
    port map (
            O => \N__28935\,
            I => \N__28913\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__28926\,
            I => \N__28910\
        );

    \I__5281\ : Span4Mux_v
    port map (
            O => \N__28921\,
            I => \N__28901\
        );

    \I__5280\ : Span4Mux_v
    port map (
            O => \N__28918\,
            I => \N__28901\
        );

    \I__5279\ : Span4Mux_h
    port map (
            O => \N__28913\,
            I => \N__28901\
        );

    \I__5278\ : Span4Mux_h
    port map (
            O => \N__28910\,
            I => \N__28901\
        );

    \I__5277\ : Span4Mux_h
    port map (
            O => \N__28901\,
            I => \N__28898\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__28898\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__28895\,
            I => \N__28891\
        );

    \I__5274\ : InMux
    port map (
            O => \N__28894\,
            I => \N__28887\
        );

    \I__5273\ : InMux
    port map (
            O => \N__28891\,
            I => \N__28884\
        );

    \I__5272\ : InMux
    port map (
            O => \N__28890\,
            I => \N__28881\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__28887\,
            I => \N__28878\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__28884\,
            I => \N__28875\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__28881\,
            I => \N__28872\
        );

    \I__5268\ : Span4Mux_h
    port map (
            O => \N__28878\,
            I => \N__28867\
        );

    \I__5267\ : Span4Mux_v
    port map (
            O => \N__28875\,
            I => \N__28867\
        );

    \I__5266\ : Span4Mux_v
    port map (
            O => \N__28872\,
            I => \N__28864\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__28867\,
            I => \il_max_comp1_D2\
        );

    \I__5264\ : Odrv4
    port map (
            O => \N__28864\,
            I => \il_max_comp1_D2\
        );

    \I__5263\ : InMux
    port map (
            O => \N__28859\,
            I => \N__28853\
        );

    \I__5262\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28845\
        );

    \I__5261\ : InMux
    port map (
            O => \N__28857\,
            I => \N__28845\
        );

    \I__5260\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28845\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__28853\,
            I => \N__28842\
        );

    \I__5258\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28839\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__28845\,
            I => \N__28835\
        );

    \I__5256\ : Span4Mux_v
    port map (
            O => \N__28842\,
            I => \N__28830\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__28839\,
            I => \N__28830\
        );

    \I__5254\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28827\
        );

    \I__5253\ : Span4Mux_h
    port map (
            O => \N__28835\,
            I => \N__28824\
        );

    \I__5252\ : Span4Mux_h
    port map (
            O => \N__28830\,
            I => \N__28821\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__28827\,
            I => state_3
        );

    \I__5250\ : Odrv4
    port map (
            O => \N__28824\,
            I => state_3
        );

    \I__5249\ : Odrv4
    port map (
            O => \N__28821\,
            I => state_3
        );

    \I__5248\ : CascadeMux
    port map (
            O => \N__28814\,
            I => \N__28810\
        );

    \I__5247\ : CascadeMux
    port map (
            O => \N__28813\,
            I => \N__28805\
        );

    \I__5246\ : InMux
    port map (
            O => \N__28810\,
            I => \N__28801\
        );

    \I__5245\ : InMux
    port map (
            O => \N__28809\,
            I => \N__28798\
        );

    \I__5244\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28794\
        );

    \I__5243\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28789\
        );

    \I__5242\ : InMux
    port map (
            O => \N__28804\,
            I => \N__28789\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__28801\,
            I => \N__28786\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__28798\,
            I => \N__28783\
        );

    \I__5239\ : InMux
    port map (
            O => \N__28797\,
            I => \N__28780\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__28794\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__28789\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5236\ : Odrv4
    port map (
            O => \N__28786\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5235\ : Odrv4
    port map (
            O => \N__28783\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__28780\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5233\ : CascadeMux
    port map (
            O => \N__28769\,
            I => \N__28766\
        );

    \I__5232\ : InMux
    port map (
            O => \N__28766\,
            I => \N__28763\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__28763\,
            I => \N__28758\
        );

    \I__5230\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28755\
        );

    \I__5229\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28752\
        );

    \I__5228\ : Span4Mux_v
    port map (
            O => \N__28758\,
            I => \N__28749\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__28755\,
            I => \N__28744\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__28752\,
            I => \N__28744\
        );

    \I__5225\ : Span4Mux_h
    port map (
            O => \N__28749\,
            I => \N__28741\
        );

    \I__5224\ : Span4Mux_v
    port map (
            O => \N__28744\,
            I => \N__28738\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__28741\,
            I => \il_min_comp1_D2\
        );

    \I__5222\ : Odrv4
    port map (
            O => \N__28738\,
            I => \il_min_comp1_D2\
        );

    \I__5221\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28729\
        );

    \I__5220\ : InMux
    port map (
            O => \N__28732\,
            I => \N__28726\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__28729\,
            I => \N__28720\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__28726\,
            I => \N__28720\
        );

    \I__5217\ : InMux
    port map (
            O => \N__28725\,
            I => \N__28717\
        );

    \I__5216\ : Span4Mux_v
    port map (
            O => \N__28720\,
            I => \N__28714\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__28717\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__5214\ : Odrv4
    port map (
            O => \N__28714\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__5213\ : InMux
    port map (
            O => \N__28709\,
            I => \N__28706\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__28706\,
            I => \N__28702\
        );

    \I__5211\ : InMux
    port map (
            O => \N__28705\,
            I => \N__28698\
        );

    \I__5210\ : Span4Mux_h
    port map (
            O => \N__28702\,
            I => \N__28695\
        );

    \I__5209\ : InMux
    port map (
            O => \N__28701\,
            I => \N__28692\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__28698\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5207\ : Odrv4
    port map (
            O => \N__28695\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__28692\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5205\ : InMux
    port map (
            O => \N__28685\,
            I => \N__28682\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__28682\,
            I => \N__28679\
        );

    \I__5203\ : Odrv12
    port map (
            O => \N__28679\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\
        );

    \I__5202\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28673\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__28673\,
            I => \N__28670\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__28670\,
            I => \N__28667\
        );

    \I__5199\ : Odrv4
    port map (
            O => \N__28667\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\
        );

    \I__5198\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28658\
        );

    \I__5197\ : InMux
    port map (
            O => \N__28663\,
            I => \N__28655\
        );

    \I__5196\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28652\
        );

    \I__5195\ : InMux
    port map (
            O => \N__28661\,
            I => \N__28649\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__28658\,
            I => \N__28646\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__28655\,
            I => \N__28641\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__28652\,
            I => \N__28641\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__28649\,
            I => \N__28637\
        );

    \I__5190\ : Span12Mux_h
    port map (
            O => \N__28646\,
            I => \N__28632\
        );

    \I__5189\ : Span12Mux_v
    port map (
            O => \N__28641\,
            I => \N__28632\
        );

    \I__5188\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28629\
        );

    \I__5187\ : Odrv4
    port map (
            O => \N__28637\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5186\ : Odrv12
    port map (
            O => \N__28632\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__28629\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5184\ : InMux
    port map (
            O => \N__28622\,
            I => \N__28619\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__28619\,
            I => \N__28616\
        );

    \I__5182\ : Span4Mux_v
    port map (
            O => \N__28616\,
            I => \N__28613\
        );

    \I__5181\ : Odrv4
    port map (
            O => \N__28613\,
            I => \current_shift_inst.un38_control_input_cry_19_c_RNOZ0\
        );

    \I__5180\ : InMux
    port map (
            O => \N__28610\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\
        );

    \I__5179\ : InMux
    port map (
            O => \N__28607\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\
        );

    \I__5178\ : InMux
    port map (
            O => \N__28604\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\
        );

    \I__5177\ : InMux
    port map (
            O => \N__28601\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_31\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__28598\,
            I => \N__28593\
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__28597\,
            I => \N__28590\
        );

    \I__5174\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28580\
        );

    \I__5173\ : InMux
    port map (
            O => \N__28593\,
            I => \N__28580\
        );

    \I__5172\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28580\
        );

    \I__5171\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28580\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__28580\,
            I => \N__28575\
        );

    \I__5169\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28572\
        );

    \I__5168\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28569\
        );

    \I__5167\ : Span4Mux_h
    port map (
            O => \N__28575\,
            I => \N__28566\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__28572\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__28569\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__28566\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__5163\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28556\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__28556\,
            I => \N__28549\
        );

    \I__5161\ : InMux
    port map (
            O => \N__28555\,
            I => \N__28540\
        );

    \I__5160\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28540\
        );

    \I__5159\ : InMux
    port map (
            O => \N__28553\,
            I => \N__28540\
        );

    \I__5158\ : InMux
    port map (
            O => \N__28552\,
            I => \N__28540\
        );

    \I__5157\ : Span4Mux_h
    port map (
            O => \N__28549\,
            I => \N__28537\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__28540\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__5155\ : Odrv4
    port map (
            O => \N__28537\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__5154\ : InMux
    port map (
            O => \N__28532\,
            I => \N__28529\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__28529\,
            I => \N__28526\
        );

    \I__5152\ : Span4Mux_v
    port map (
            O => \N__28526\,
            I => \N__28523\
        );

    \I__5151\ : Odrv4
    port map (
            O => \N__28523\,
            I => \phase_controller_inst1.stoper_tr.N_45\
        );

    \I__5150\ : InMux
    port map (
            O => \N__28520\,
            I => \N__28516\
        );

    \I__5149\ : InMux
    port map (
            O => \N__28519\,
            I => \N__28513\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__28516\,
            I => \N__28510\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__28513\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5146\ : Odrv12
    port map (
            O => \N__28510\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5145\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28502\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__28502\,
            I => \N__28499\
        );

    \I__5143\ : Odrv12
    port map (
            O => \N__28499\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\
        );

    \I__5142\ : InMux
    port map (
            O => \N__28496\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\
        );

    \I__5141\ : InMux
    port map (
            O => \N__28493\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\
        );

    \I__5140\ : InMux
    port map (
            O => \N__28490\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\
        );

    \I__5139\ : InMux
    port map (
            O => \N__28487\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\
        );

    \I__5138\ : InMux
    port map (
            O => \N__28484\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\
        );

    \I__5137\ : InMux
    port map (
            O => \N__28481\,
            I => \bfn_13_14_0_\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__28478\,
            I => \N__28475\
        );

    \I__5135\ : InMux
    port map (
            O => \N__28475\,
            I => \N__28472\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__28472\,
            I => \N__28469\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__28469\,
            I => \N__28466\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__28466\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\
        );

    \I__5131\ : InMux
    port map (
            O => \N__28463\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\
        );

    \I__5130\ : InMux
    port map (
            O => \N__28460\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\
        );

    \I__5129\ : InMux
    port map (
            O => \N__28457\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\
        );

    \I__5128\ : InMux
    port map (
            O => \N__28454\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\
        );

    \I__5127\ : InMux
    port map (
            O => \N__28451\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\
        );

    \I__5126\ : InMux
    port map (
            O => \N__28448\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\
        );

    \I__5125\ : InMux
    port map (
            O => \N__28445\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\
        );

    \I__5124\ : InMux
    port map (
            O => \N__28442\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\
        );

    \I__5123\ : InMux
    port map (
            O => \N__28439\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\
        );

    \I__5122\ : InMux
    port map (
            O => \N__28436\,
            I => \bfn_13_13_0_\
        );

    \I__5121\ : InMux
    port map (
            O => \N__28433\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\
        );

    \I__5120\ : InMux
    port map (
            O => \N__28430\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\
        );

    \I__5119\ : InMux
    port map (
            O => \N__28427\,
            I => \N__28424\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__28424\,
            I => \N__28420\
        );

    \I__5117\ : InMux
    port map (
            O => \N__28423\,
            I => \N__28417\
        );

    \I__5116\ : Span4Mux_h
    port map (
            O => \N__28420\,
            I => \N__28414\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__28417\,
            I => \N__28411\
        );

    \I__5114\ : Odrv4
    port map (
            O => \N__28414\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__28411\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__5112\ : InMux
    port map (
            O => \N__28406\,
            I => \N__28403\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__28403\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\
        );

    \I__5110\ : InMux
    port map (
            O => \N__28400\,
            I => \N__28397\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__28397\,
            I => \N__28394\
        );

    \I__5108\ : Span4Mux_h
    port map (
            O => \N__28394\,
            I => \N__28390\
        );

    \I__5107\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28387\
        );

    \I__5106\ : Odrv4
    port map (
            O => \N__28390\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__28387\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__5104\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28379\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__28379\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\
        );

    \I__5102\ : InMux
    port map (
            O => \N__28376\,
            I => \N__28373\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__28373\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__28370\,
            I => \N__28367\
        );

    \I__5099\ : InMux
    port map (
            O => \N__28367\,
            I => \N__28364\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__28364\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_4\
        );

    \I__5097\ : InMux
    port map (
            O => \N__28361\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\
        );

    \I__5096\ : InMux
    port map (
            O => \N__28358\,
            I => \N__28355\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__28355\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\
        );

    \I__5094\ : CascadeMux
    port map (
            O => \N__28352\,
            I => \N__28349\
        );

    \I__5093\ : InMux
    port map (
            O => \N__28349\,
            I => \N__28346\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__28346\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_5\
        );

    \I__5091\ : InMux
    port map (
            O => \N__28343\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\
        );

    \I__5090\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28337\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__28337\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\
        );

    \I__5088\ : InMux
    port map (
            O => \N__28334\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\
        );

    \I__5087\ : InMux
    port map (
            O => \N__28331\,
            I => \N__28328\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__28328\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\
        );

    \I__5085\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28322\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__28322\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_7\
        );

    \I__5083\ : InMux
    port map (
            O => \N__28319\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\
        );

    \I__5082\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28313\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__28313\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\
        );

    \I__5080\ : InMux
    port map (
            O => \N__28310\,
            I => \bfn_13_12_0_\
        );

    \I__5079\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28304\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__28304\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\
        );

    \I__5077\ : InMux
    port map (
            O => \N__28301\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\
        );

    \I__5076\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28295\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__28295\,
            I => \N__28292\
        );

    \I__5074\ : Span4Mux_h
    port map (
            O => \N__28292\,
            I => \N__28287\
        );

    \I__5073\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28282\
        );

    \I__5072\ : InMux
    port map (
            O => \N__28290\,
            I => \N__28282\
        );

    \I__5071\ : Odrv4
    port map (
            O => \N__28287\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__28282\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5069\ : InMux
    port map (
            O => \N__28277\,
            I => \N__28274\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__28274\,
            I => \N__28271\
        );

    \I__5067\ : Span4Mux_h
    port map (
            O => \N__28271\,
            I => \N__28266\
        );

    \I__5066\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28261\
        );

    \I__5065\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28261\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__28266\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__28261\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__5062\ : InMux
    port map (
            O => \N__28256\,
            I => \N__28253\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__28253\,
            I => \N__28249\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28252\,
            I => \N__28246\
        );

    \I__5059\ : Span4Mux_h
    port map (
            O => \N__28249\,
            I => \N__28241\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__28246\,
            I => \N__28241\
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__28241\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__5056\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28235\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__28235\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\
        );

    \I__5054\ : InMux
    port map (
            O => \N__28232\,
            I => \N__28228\
        );

    \I__5053\ : InMux
    port map (
            O => \N__28231\,
            I => \N__28225\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__28228\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__28225\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__5050\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28217\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__28217\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\
        );

    \I__5048\ : InMux
    port map (
            O => \N__28214\,
            I => \N__28211\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__28211\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\
        );

    \I__5046\ : InMux
    port map (
            O => \N__28208\,
            I => \N__28205\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__28205\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__5044\ : InMux
    port map (
            O => \N__28202\,
            I => \N__28199\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__28199\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__5042\ : CascadeMux
    port map (
            O => \N__28196\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19_cascade_\
        );

    \I__5041\ : CascadeMux
    port map (
            O => \N__28193\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\
        );

    \I__5040\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28187\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__28187\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\
        );

    \I__5038\ : InMux
    port map (
            O => \N__28184\,
            I => \N__28181\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__28181\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16\
        );

    \I__5036\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28175\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__28175\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\
        );

    \I__5034\ : InMux
    port map (
            O => \N__28172\,
            I => \N__28169\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__28169\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__5032\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28162\
        );

    \I__5031\ : InMux
    port map (
            O => \N__28165\,
            I => \N__28159\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__28162\,
            I => \current_shift_inst.PI_CTRL.N_74_21\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__28159\,
            I => \current_shift_inst.PI_CTRL.N_74_21\
        );

    \I__5028\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28151\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__28151\,
            I => \N__28148\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__28148\,
            I => \N__28144\
        );

    \I__5025\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28141\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__28144\,
            I => \current_shift_inst.PI_CTRL.N_72\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__28141\,
            I => \current_shift_inst.PI_CTRL.N_72\
        );

    \I__5022\ : InMux
    port map (
            O => \N__28136\,
            I => \N__28133\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__28133\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__5020\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28120\
        );

    \I__5019\ : InMux
    port map (
            O => \N__28129\,
            I => \N__28120\
        );

    \I__5018\ : InMux
    port map (
            O => \N__28128\,
            I => \N__28120\
        );

    \I__5017\ : InMux
    port map (
            O => \N__28127\,
            I => \N__28117\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__28120\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__28117\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__5014\ : InMux
    port map (
            O => \N__28112\,
            I => \N__28106\
        );

    \I__5013\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28099\
        );

    \I__5012\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28099\
        );

    \I__5011\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28099\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__28106\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__28099\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__28094\,
            I => \N__28091\
        );

    \I__5007\ : InMux
    port map (
            O => \N__28091\,
            I => \N__28083\
        );

    \I__5006\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28083\
        );

    \I__5005\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28078\
        );

    \I__5004\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28078\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__28083\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__28078\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__5001\ : IoInMux
    port map (
            O => \N__28073\,
            I => \N__28070\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__28070\,
            I => \N__28067\
        );

    \I__4999\ : IoSpan4Mux
    port map (
            O => \N__28067\,
            I => \N__28064\
        );

    \I__4998\ : Span4Mux_s0_v
    port map (
            O => \N__28064\,
            I => \N__28061\
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__28061\,
            I => \pll_inst.red_c_i\
        );

    \I__4996\ : CascadeMux
    port map (
            O => \N__28058\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18_cascade_\
        );

    \I__4995\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28052\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__28052\,
            I => \current_shift_inst.PI_CTRL.N_62\
        );

    \I__4993\ : CascadeMux
    port map (
            O => \N__28049\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_\
        );

    \I__4992\ : InMux
    port map (
            O => \N__28046\,
            I => \N__28040\
        );

    \I__4991\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28040\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__28040\,
            I => \current_shift_inst.un38_control_input_axb_30\
        );

    \I__4989\ : InMux
    port map (
            O => \N__28037\,
            I => \N__28033\
        );

    \I__4988\ : InMux
    port map (
            O => \N__28036\,
            I => \N__28030\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__28033\,
            I => \N__28027\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__28030\,
            I => \N__28024\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__28027\,
            I => \phase_controller_inst2.time_passed_RNI9M3O\
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__28024\,
            I => \phase_controller_inst2.time_passed_RNI9M3O\
        );

    \I__4983\ : InMux
    port map (
            O => \N__28019\,
            I => \N__28016\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__28016\,
            I => \N__28012\
        );

    \I__4981\ : InMux
    port map (
            O => \N__28015\,
            I => \N__28006\
        );

    \I__4980\ : Span4Mux_h
    port map (
            O => \N__28012\,
            I => \N__28003\
        );

    \I__4979\ : InMux
    port map (
            O => \N__28011\,
            I => \N__28000\
        );

    \I__4978\ : InMux
    port map (
            O => \N__28010\,
            I => \N__27995\
        );

    \I__4977\ : InMux
    port map (
            O => \N__28009\,
            I => \N__27995\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__28006\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4975\ : Odrv4
    port map (
            O => \N__28003\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__28000\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__27995\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4972\ : IoInMux
    port map (
            O => \N__27986\,
            I => \N__27983\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__27983\,
            I => \N__27980\
        );

    \I__4970\ : Span4Mux_s3_v
    port map (
            O => \N__27980\,
            I => \N__27977\
        );

    \I__4969\ : Span4Mux_h
    port map (
            O => \N__27977\,
            I => \N__27974\
        );

    \I__4968\ : Span4Mux_v
    port map (
            O => \N__27974\,
            I => \N__27970\
        );

    \I__4967\ : InMux
    port map (
            O => \N__27973\,
            I => \N__27967\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__27970\,
            I => \T01_c\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__27967\,
            I => \T01_c\
        );

    \I__4964\ : IoInMux
    port map (
            O => \N__27962\,
            I => \N__27959\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__27959\,
            I => \N__27956\
        );

    \I__4962\ : Span4Mux_s1_v
    port map (
            O => \N__27956\,
            I => \N__27953\
        );

    \I__4961\ : Span4Mux_v
    port map (
            O => \N__27953\,
            I => \N__27948\
        );

    \I__4960\ : InMux
    port map (
            O => \N__27952\,
            I => \N__27943\
        );

    \I__4959\ : InMux
    port map (
            O => \N__27951\,
            I => \N__27943\
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__27948\,
            I => s1_phy_c
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__27943\,
            I => s1_phy_c
        );

    \I__4956\ : CascadeMux
    port map (
            O => \N__27938\,
            I => \N__27933\
        );

    \I__4955\ : InMux
    port map (
            O => \N__27937\,
            I => \N__27930\
        );

    \I__4954\ : InMux
    port map (
            O => \N__27936\,
            I => \N__27926\
        );

    \I__4953\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27923\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__27930\,
            I => \N__27920\
        );

    \I__4951\ : InMux
    port map (
            O => \N__27929\,
            I => \N__27917\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__27926\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__27923\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__4948\ : Odrv4
    port map (
            O => \N__27920\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__27917\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__4946\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27902\
        );

    \I__4945\ : InMux
    port map (
            O => \N__27907\,
            I => \N__27899\
        );

    \I__4944\ : InMux
    port map (
            O => \N__27906\,
            I => \N__27896\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__27905\,
            I => \N__27892\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__27902\,
            I => \N__27888\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__27899\,
            I => \N__27885\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__27896\,
            I => \N__27882\
        );

    \I__4939\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27879\
        );

    \I__4938\ : InMux
    port map (
            O => \N__27892\,
            I => \N__27876\
        );

    \I__4937\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27873\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__27888\,
            I => \N__27868\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__27885\,
            I => \N__27868\
        );

    \I__4934\ : Span4Mux_h
    port map (
            O => \N__27882\,
            I => \N__27863\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__27879\,
            I => \N__27863\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__27876\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__27873\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__27868\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__27863\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4928\ : IoInMux
    port map (
            O => \N__27854\,
            I => \N__27851\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__27851\,
            I => \N__27848\
        );

    \I__4926\ : Span4Mux_s2_v
    port map (
            O => \N__27848\,
            I => \N__27845\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__27845\,
            I => \N__27841\
        );

    \I__4924\ : InMux
    port map (
            O => \N__27844\,
            I => \N__27838\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__27841\,
            I => \T45_c\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__27838\,
            I => \T45_c\
        );

    \I__4921\ : IoInMux
    port map (
            O => \N__27833\,
            I => \N__27830\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__27830\,
            I => \N__27827\
        );

    \I__4919\ : Span4Mux_s1_v
    port map (
            O => \N__27827\,
            I => \N__27824\
        );

    \I__4918\ : Odrv4
    port map (
            O => \N__27824\,
            I => \current_shift_inst.timer_s1.N_166_i\
        );

    \I__4917\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27818\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__27818\,
            I => \current_shift_inst.control_input_1_axb_3\
        );

    \I__4915\ : InMux
    port map (
            O => \N__27815\,
            I => \bfn_12_21_0_\
        );

    \I__4914\ : InMux
    port map (
            O => \N__27812\,
            I => \N__27809\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__27809\,
            I => \current_shift_inst.control_input_1_axb_4\
        );

    \I__4912\ : InMux
    port map (
            O => \N__27806\,
            I => \current_shift_inst.un38_control_input_cry_23\
        );

    \I__4911\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27800\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__27800\,
            I => \current_shift_inst.control_input_1_axb_5\
        );

    \I__4909\ : InMux
    port map (
            O => \N__27797\,
            I => \current_shift_inst.un38_control_input_cry_24\
        );

    \I__4908\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27791\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__27791\,
            I => \current_shift_inst.control_input_1_axb_6\
        );

    \I__4906\ : InMux
    port map (
            O => \N__27788\,
            I => \current_shift_inst.un38_control_input_cry_25\
        );

    \I__4905\ : InMux
    port map (
            O => \N__27785\,
            I => \N__27782\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__27782\,
            I => \N__27779\
        );

    \I__4903\ : Span4Mux_v
    port map (
            O => \N__27779\,
            I => \N__27776\
        );

    \I__4902\ : Odrv4
    port map (
            O => \N__27776\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__4901\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27770\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__27770\,
            I => \current_shift_inst.control_input_1_axb_7\
        );

    \I__4899\ : InMux
    port map (
            O => \N__27767\,
            I => \current_shift_inst.un38_control_input_cry_26\
        );

    \I__4898\ : InMux
    port map (
            O => \N__27764\,
            I => \N__27761\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__27761\,
            I => \current_shift_inst.control_input_1_axb_8\
        );

    \I__4896\ : InMux
    port map (
            O => \N__27758\,
            I => \current_shift_inst.un38_control_input_cry_27\
        );

    \I__4895\ : InMux
    port map (
            O => \N__27755\,
            I => \N__27752\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__27752\,
            I => \current_shift_inst.control_input_1_axb_9\
        );

    \I__4893\ : InMux
    port map (
            O => \N__27749\,
            I => \current_shift_inst.un38_control_input_cry_28\
        );

    \I__4892\ : InMux
    port map (
            O => \N__27746\,
            I => \current_shift_inst.un38_control_input_cry_29\
        );

    \I__4891\ : CascadeMux
    port map (
            O => \N__27743\,
            I => \N__27740\
        );

    \I__4890\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27736\
        );

    \I__4889\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27733\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__27736\,
            I => \current_shift_inst.un38_control_input_cry_29_THRU_CO\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__27733\,
            I => \current_shift_inst.un38_control_input_cry_29_THRU_CO\
        );

    \I__4886\ : InMux
    port map (
            O => \N__27728\,
            I => \N__27725\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__27725\,
            I => \current_shift_inst.control_input_1_axb_0\
        );

    \I__4884\ : InMux
    port map (
            O => \N__27722\,
            I => \current_shift_inst.un38_control_input_cry_19\
        );

    \I__4883\ : InMux
    port map (
            O => \N__27719\,
            I => \N__27716\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__27716\,
            I => \current_shift_inst.control_input_1_axb_1\
        );

    \I__4881\ : InMux
    port map (
            O => \N__27713\,
            I => \current_shift_inst.un38_control_input_cry_20\
        );

    \I__4880\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27707\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__27707\,
            I => \current_shift_inst.control_input_1_axb_2\
        );

    \I__4878\ : InMux
    port map (
            O => \N__27704\,
            I => \current_shift_inst.un38_control_input_cry_21\
        );

    \I__4877\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27698\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__27698\,
            I => \N__27695\
        );

    \I__4875\ : Odrv12
    port map (
            O => \N__27695\,
            I => \current_shift_inst.un38_control_input_cry_7_c_RNOZ0\
        );

    \I__4874\ : InMux
    port map (
            O => \N__27692\,
            I => \N__27689\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__27689\,
            I => \current_shift_inst.un38_control_input_cry_3_c_RNOZ0\
        );

    \I__4872\ : InMux
    port map (
            O => \N__27686\,
            I => \N__27683\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__27683\,
            I => \current_shift_inst.un38_control_input_cry_4_c_RNOZ0\
        );

    \I__4870\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27676\
        );

    \I__4869\ : InMux
    port map (
            O => \N__27679\,
            I => \N__27673\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__27676\,
            I => \N__27670\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__27673\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4866\ : Odrv4
    port map (
            O => \N__27670\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4865\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27662\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__27662\,
            I => \N__27659\
        );

    \I__4863\ : Span4Mux_h
    port map (
            O => \N__27659\,
            I => \N__27656\
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__27656\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__4861\ : CascadeMux
    port map (
            O => \N__27653\,
            I => \N__27650\
        );

    \I__4860\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27647\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__27647\,
            I => \N__27644\
        );

    \I__4858\ : Odrv4
    port map (
            O => \N__27644\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__4857\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27638\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__27638\,
            I => \N__27635\
        );

    \I__4855\ : Span4Mux_h
    port map (
            O => \N__27635\,
            I => \N__27632\
        );

    \I__4854\ : Odrv4
    port map (
            O => \N__27632\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__4853\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27625\
        );

    \I__4852\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27622\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__27625\,
            I => \N__27619\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__27622\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__27619\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__27614\,
            I => \N__27611\
        );

    \I__4847\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27608\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__27608\,
            I => \N__27605\
        );

    \I__4845\ : Odrv4
    port map (
            O => \N__27605\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__4844\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27598\
        );

    \I__4843\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27595\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__27598\,
            I => \N__27592\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__27595\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__27592\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4839\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27584\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__27584\,
            I => \N__27581\
        );

    \I__4837\ : Span4Mux_v
    port map (
            O => \N__27581\,
            I => \N__27578\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__27578\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__4835\ : CascadeMux
    port map (
            O => \N__27575\,
            I => \N__27572\
        );

    \I__4834\ : InMux
    port map (
            O => \N__27572\,
            I => \N__27569\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__27569\,
            I => \N__27566\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__27566\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\
        );

    \I__4831\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27559\
        );

    \I__4830\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27556\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__27559\,
            I => \N__27553\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__27556\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__27553\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4826\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27545\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__4824\ : Span4Mux_h
    port map (
            O => \N__27542\,
            I => \N__27539\
        );

    \I__4823\ : Odrv4
    port map (
            O => \N__27539\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__4822\ : CascadeMux
    port map (
            O => \N__27536\,
            I => \N__27533\
        );

    \I__4821\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27530\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__27530\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\
        );

    \I__4819\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27523\
        );

    \I__4818\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27520\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__27523\,
            I => \N__27517\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__27520\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__27517\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4814\ : InMux
    port map (
            O => \N__27512\,
            I => \N__27509\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__27509\,
            I => \N__27506\
        );

    \I__4812\ : Span4Mux_v
    port map (
            O => \N__27506\,
            I => \N__27503\
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__27503\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__4810\ : CascadeMux
    port map (
            O => \N__27500\,
            I => \N__27497\
        );

    \I__4809\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27494\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__27494\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\
        );

    \I__4807\ : InMux
    port map (
            O => \N__27491\,
            I => \N__27488\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__27488\,
            I => \N__27485\
        );

    \I__4805\ : Span4Mux_v
    port map (
            O => \N__27485\,
            I => \N__27482\
        );

    \I__4804\ : Odrv4
    port map (
            O => \N__27482\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__4803\ : InMux
    port map (
            O => \N__27479\,
            I => \N__27475\
        );

    \I__4802\ : InMux
    port map (
            O => \N__27478\,
            I => \N__27472\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__27475\,
            I => \N__27469\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__27472\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4799\ : Odrv4
    port map (
            O => \N__27469\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4798\ : CascadeMux
    port map (
            O => \N__27464\,
            I => \N__27461\
        );

    \I__4797\ : InMux
    port map (
            O => \N__27461\,
            I => \N__27458\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__27458\,
            I => \N__27455\
        );

    \I__4795\ : Odrv4
    port map (
            O => \N__27455\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\
        );

    \I__4794\ : InMux
    port map (
            O => \N__27452\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__4793\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27446\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__27446\,
            I => \N__27442\
        );

    \I__4791\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27439\
        );

    \I__4790\ : Span4Mux_h
    port map (
            O => \N__27442\,
            I => \N__27436\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__27439\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__4788\ : Odrv4
    port map (
            O => \N__27436\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__4787\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27428\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__27428\,
            I => \N__27425\
        );

    \I__4785\ : Span4Mux_v
    port map (
            O => \N__27425\,
            I => \N__27422\
        );

    \I__4784\ : Odrv4
    port map (
            O => \N__27422\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__4783\ : CascadeMux
    port map (
            O => \N__27419\,
            I => \N__27416\
        );

    \I__4782\ : InMux
    port map (
            O => \N__27416\,
            I => \N__27413\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__27413\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__4780\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27407\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__27407\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__4778\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27400\
        );

    \I__4777\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27397\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__27400\,
            I => \N__27394\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__27397\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__27394\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__27389\,
            I => \N__27386\
        );

    \I__4772\ : InMux
    port map (
            O => \N__27386\,
            I => \N__27383\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__27383\,
            I => \N__27380\
        );

    \I__4770\ : Odrv12
    port map (
            O => \N__27380\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__4769\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27373\
        );

    \I__4768\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27370\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__27373\,
            I => \N__27367\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__27370\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__27367\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__4764\ : InMux
    port map (
            O => \N__27362\,
            I => \N__27359\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__27359\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__4762\ : CascadeMux
    port map (
            O => \N__27356\,
            I => \N__27353\
        );

    \I__4761\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27350\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__27350\,
            I => \N__27347\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__27347\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__4758\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27341\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__27341\,
            I => \N__27338\
        );

    \I__4756\ : Span12Mux_h
    port map (
            O => \N__27338\,
            I => \N__27335\
        );

    \I__4755\ : Odrv12
    port map (
            O => \N__27335\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__4754\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27329\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__27329\,
            I => \N__27326\
        );

    \I__4752\ : Span4Mux_h
    port map (
            O => \N__27326\,
            I => \N__27322\
        );

    \I__4751\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27319\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__27322\,
            I => \N__27316\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__27319\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4748\ : Odrv4
    port map (
            O => \N__27316\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__27311\,
            I => \N__27308\
        );

    \I__4746\ : InMux
    port map (
            O => \N__27308\,
            I => \N__27305\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__27305\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__4744\ : InMux
    port map (
            O => \N__27302\,
            I => \N__27299\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__27299\,
            I => \N__27296\
        );

    \I__4742\ : Span4Mux_h
    port map (
            O => \N__27296\,
            I => \N__27293\
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__27293\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__4740\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27286\
        );

    \I__4739\ : InMux
    port map (
            O => \N__27289\,
            I => \N__27283\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__27286\,
            I => \N__27280\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__27283\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4736\ : Odrv4
    port map (
            O => \N__27280\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__27275\,
            I => \N__27272\
        );

    \I__4734\ : InMux
    port map (
            O => \N__27272\,
            I => \N__27269\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__27269\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__4732\ : InMux
    port map (
            O => \N__27266\,
            I => \N__27263\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__27263\,
            I => \N__27259\
        );

    \I__4730\ : InMux
    port map (
            O => \N__27262\,
            I => \N__27256\
        );

    \I__4729\ : Span4Mux_v
    port map (
            O => \N__27259\,
            I => \N__27253\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__27256\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4727\ : Odrv4
    port map (
            O => \N__27253\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4726\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27245\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__27245\,
            I => \N__27242\
        );

    \I__4724\ : Span4Mux_h
    port map (
            O => \N__27242\,
            I => \N__27239\
        );

    \I__4723\ : Odrv4
    port map (
            O => \N__27239\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__4722\ : CascadeMux
    port map (
            O => \N__27236\,
            I => \N__27233\
        );

    \I__4721\ : InMux
    port map (
            O => \N__27233\,
            I => \N__27230\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__27230\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__4719\ : InMux
    port map (
            O => \N__27227\,
            I => \N__27224\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__27224\,
            I => \N__27221\
        );

    \I__4717\ : Span4Mux_h
    port map (
            O => \N__27221\,
            I => \N__27218\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__27218\,
            I => \N__27215\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__27215\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__4714\ : InMux
    port map (
            O => \N__27212\,
            I => \N__27208\
        );

    \I__4713\ : InMux
    port map (
            O => \N__27211\,
            I => \N__27205\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__27208\,
            I => \N__27202\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__27205\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__27202\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4709\ : CascadeMux
    port map (
            O => \N__27197\,
            I => \N__27194\
        );

    \I__4708\ : InMux
    port map (
            O => \N__27194\,
            I => \N__27191\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__27191\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__4706\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27184\
        );

    \I__4705\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27181\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__27184\,
            I => \N__27178\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__27181\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4702\ : Odrv4
    port map (
            O => \N__27178\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4701\ : InMux
    port map (
            O => \N__27173\,
            I => \N__27170\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__27170\,
            I => \N__27167\
        );

    \I__4699\ : Span4Mux_v
    port map (
            O => \N__27167\,
            I => \N__27164\
        );

    \I__4698\ : Span4Mux_h
    port map (
            O => \N__27164\,
            I => \N__27161\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__27161\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__27158\,
            I => \N__27155\
        );

    \I__4695\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27152\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__27152\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__4693\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27146\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__27146\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__4691\ : CascadeMux
    port map (
            O => \N__27143\,
            I => \N__27140\
        );

    \I__4690\ : InMux
    port map (
            O => \N__27140\,
            I => \N__27137\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__27137\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__4688\ : CascadeMux
    port map (
            O => \N__27134\,
            I => \N__27131\
        );

    \I__4687\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27128\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__27128\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__4685\ : InMux
    port map (
            O => \N__27125\,
            I => \N__27121\
        );

    \I__4684\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27118\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__27121\,
            I => \N__27115\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__27118\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4681\ : Odrv4
    port map (
            O => \N__27115\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4680\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27107\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__27107\,
            I => \N__27104\
        );

    \I__4678\ : Odrv4
    port map (
            O => \N__27104\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__27101\,
            I => \N__27097\
        );

    \I__4676\ : InMux
    port map (
            O => \N__27100\,
            I => \N__27094\
        );

    \I__4675\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27091\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__27094\,
            I => \N__27088\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__27091\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__27088\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__27083\,
            I => \N__27080\
        );

    \I__4670\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27077\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__27077\,
            I => \N__27074\
        );

    \I__4668\ : Span4Mux_h
    port map (
            O => \N__27074\,
            I => \N__27071\
        );

    \I__4667\ : Odrv4
    port map (
            O => \N__27071\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__4666\ : InMux
    port map (
            O => \N__27068\,
            I => \N__27065\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__27065\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__4664\ : InMux
    port map (
            O => \N__27062\,
            I => \N__27059\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__27059\,
            I => \N__27056\
        );

    \I__4662\ : Span4Mux_h
    port map (
            O => \N__27056\,
            I => \N__27053\
        );

    \I__4661\ : Odrv4
    port map (
            O => \N__27053\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__4660\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27046\
        );

    \I__4659\ : InMux
    port map (
            O => \N__27049\,
            I => \N__27043\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__27046\,
            I => \N__27040\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__27043\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__27040\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__27035\,
            I => \N__27032\
        );

    \I__4654\ : InMux
    port map (
            O => \N__27032\,
            I => \N__27029\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__27029\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__4652\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27022\
        );

    \I__4651\ : InMux
    port map (
            O => \N__27025\,
            I => \N__27019\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__27022\,
            I => \N__27016\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__27019\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__27016\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__4647\ : InMux
    port map (
            O => \N__27011\,
            I => \N__27008\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__27008\,
            I => \N__27005\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__27005\,
            I => \N__27002\
        );

    \I__4644\ : Odrv4
    port map (
            O => \N__27002\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__4643\ : CascadeMux
    port map (
            O => \N__26999\,
            I => \N__26996\
        );

    \I__4642\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26993\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__26993\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__4640\ : InMux
    port map (
            O => \N__26990\,
            I => \N__26987\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__26987\,
            I => \N__26984\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__26984\,
            I => \N__26981\
        );

    \I__4637\ : Span4Mux_v
    port map (
            O => \N__26981\,
            I => \N__26978\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__26978\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__4635\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26972\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__26972\,
            I => \N__26969\
        );

    \I__4633\ : Odrv4
    port map (
            O => \N__26969\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__4632\ : InMux
    port map (
            O => \N__26966\,
            I => \N__26963\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__26963\,
            I => \N__26960\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__26960\,
            I => \N__26957\
        );

    \I__4629\ : Span4Mux_v
    port map (
            O => \N__26957\,
            I => \N__26954\
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__26954\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__4627\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26948\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__26948\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__4625\ : InMux
    port map (
            O => \N__26945\,
            I => \N__26942\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__26942\,
            I => \N__26939\
        );

    \I__4623\ : Span4Mux_v
    port map (
            O => \N__26939\,
            I => \N__26936\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__26936\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__4621\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26930\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__26930\,
            I => \N__26927\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__26927\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__4618\ : InMux
    port map (
            O => \N__26924\,
            I => \N__26921\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__26921\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHEZ0\
        );

    \I__4616\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26915\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__26915\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__4614\ : InMux
    port map (
            O => \N__26912\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__4613\ : InMux
    port map (
            O => \N__26909\,
            I => \N__26906\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__26906\,
            I => \N__26903\
        );

    \I__4611\ : Span4Mux_h
    port map (
            O => \N__26903\,
            I => \N__26898\
        );

    \I__4610\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26893\
        );

    \I__4609\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26893\
        );

    \I__4608\ : Odrv4
    port map (
            O => \N__26898\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__26893\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__4606\ : InMux
    port map (
            O => \N__26888\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__4605\ : InMux
    port map (
            O => \N__26885\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__4604\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26879\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__26879\,
            I => \N__26876\
        );

    \I__4602\ : Span12Mux_v
    port map (
            O => \N__26876\,
            I => \N__26873\
        );

    \I__4601\ : Odrv12
    port map (
            O => \N__26873\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__4600\ : InMux
    port map (
            O => \N__26870\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__4599\ : InMux
    port map (
            O => \N__26867\,
            I => \bfn_12_12_0_\
        );

    \I__4598\ : InMux
    port map (
            O => \N__26864\,
            I => \N__26861\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__26861\,
            I => \N__26858\
        );

    \I__4596\ : Span4Mux_v
    port map (
            O => \N__26858\,
            I => \N__26855\
        );

    \I__4595\ : Span4Mux_v
    port map (
            O => \N__26855\,
            I => \N__26852\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__26852\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__4593\ : InMux
    port map (
            O => \N__26849\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__4592\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26843\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__26843\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__4590\ : InMux
    port map (
            O => \N__26840\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__4589\ : InMux
    port map (
            O => \N__26837\,
            I => \N__26834\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__26834\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__4587\ : InMux
    port map (
            O => \N__26831\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__4586\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26825\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__26825\,
            I => \N__26821\
        );

    \I__4584\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26818\
        );

    \I__4583\ : Span4Mux_h
    port map (
            O => \N__26821\,
            I => \N__26815\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__26818\,
            I => \N__26812\
        );

    \I__4581\ : Sp12to4
    port map (
            O => \N__26815\,
            I => \N__26807\
        );

    \I__4580\ : Span12Mux_v
    port map (
            O => \N__26812\,
            I => \N__26807\
        );

    \I__4579\ : Odrv12
    port map (
            O => \N__26807\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__4578\ : InMux
    port map (
            O => \N__26804\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__4577\ : InMux
    port map (
            O => \N__26801\,
            I => \N__26798\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__26798\,
            I => \N__26794\
        );

    \I__4575\ : InMux
    port map (
            O => \N__26797\,
            I => \N__26791\
        );

    \I__4574\ : Span4Mux_v
    port map (
            O => \N__26794\,
            I => \N__26788\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__26791\,
            I => \N__26785\
        );

    \I__4572\ : Span4Mux_v
    port map (
            O => \N__26788\,
            I => \N__26782\
        );

    \I__4571\ : Odrv12
    port map (
            O => \N__26785\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__26782\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__4569\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__26774\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__4567\ : InMux
    port map (
            O => \N__26771\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__4566\ : InMux
    port map (
            O => \N__26768\,
            I => \N__26765\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__26765\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__4564\ : InMux
    port map (
            O => \N__26762\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__4563\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26756\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__26756\,
            I => \N__26753\
        );

    \I__4561\ : Span4Mux_v
    port map (
            O => \N__26753\,
            I => \N__26750\
        );

    \I__4560\ : Odrv4
    port map (
            O => \N__26750\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__4559\ : InMux
    port map (
            O => \N__26747\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__26744\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_\
        );

    \I__4557\ : InMux
    port map (
            O => \N__26741\,
            I => \N__26738\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__26738\,
            I => \N__26735\
        );

    \I__4555\ : Odrv4
    port map (
            O => \N__26735\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__26732\,
            I => \current_shift_inst.PI_CTRL.N_74_16_cascade_\
        );

    \I__4553\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26726\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__26726\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__4551\ : InMux
    port map (
            O => \N__26723\,
            I => \N__26720\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__26720\,
            I => \N__26716\
        );

    \I__4549\ : InMux
    port map (
            O => \N__26719\,
            I => \N__26713\
        );

    \I__4548\ : Span4Mux_s1_v
    port map (
            O => \N__26716\,
            I => \N__26708\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__26713\,
            I => \N__26708\
        );

    \I__4546\ : Span4Mux_v
    port map (
            O => \N__26708\,
            I => \N__26705\
        );

    \I__4545\ : Span4Mux_h
    port map (
            O => \N__26705\,
            I => \N__26702\
        );

    \I__4544\ : Sp12to4
    port map (
            O => \N__26702\,
            I => \N__26697\
        );

    \I__4543\ : InMux
    port map (
            O => \N__26701\,
            I => \N__26694\
        );

    \I__4542\ : InMux
    port map (
            O => \N__26700\,
            I => \N__26691\
        );

    \I__4541\ : Span12Mux_v
    port map (
            O => \N__26697\,
            I => \N__26688\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__26694\,
            I => \N__26683\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__26691\,
            I => \N__26683\
        );

    \I__4538\ : Span12Mux_v
    port map (
            O => \N__26688\,
            I => \N__26680\
        );

    \I__4537\ : Span12Mux_h
    port map (
            O => \N__26683\,
            I => \N__26677\
        );

    \I__4536\ : Span12Mux_h
    port map (
            O => \N__26680\,
            I => \N__26674\
        );

    \I__4535\ : Span12Mux_v
    port map (
            O => \N__26677\,
            I => \N__26671\
        );

    \I__4534\ : Odrv12
    port map (
            O => \N__26674\,
            I => start_stop_c
        );

    \I__4533\ : Odrv12
    port map (
            O => \N__26671\,
            I => start_stop_c
        );

    \I__4532\ : InMux
    port map (
            O => \N__26666\,
            I => \N__26660\
        );

    \I__4531\ : InMux
    port map (
            O => \N__26665\,
            I => \N__26657\
        );

    \I__4530\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26652\
        );

    \I__4529\ : InMux
    port map (
            O => \N__26663\,
            I => \N__26652\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__26660\,
            I => \N__26647\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__26657\,
            I => \N__26642\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__26652\,
            I => \N__26642\
        );

    \I__4525\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26639\
        );

    \I__4524\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26636\
        );

    \I__4523\ : Odrv12
    port map (
            O => \N__26647\,
            I => phase_controller_inst1_state_4
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__26642\,
            I => phase_controller_inst1_state_4
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__26639\,
            I => phase_controller_inst1_state_4
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__26636\,
            I => phase_controller_inst1_state_4
        );

    \I__4519\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26624\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__26624\,
            I => \N__26619\
        );

    \I__4517\ : InMux
    port map (
            O => \N__26623\,
            I => \N__26614\
        );

    \I__4516\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26614\
        );

    \I__4515\ : Span4Mux_h
    port map (
            O => \N__26619\,
            I => \N__26611\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__26614\,
            I => \N__26608\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__26611\,
            I => \il_min_comp2_D2\
        );

    \I__4512\ : Odrv12
    port map (
            O => \N__26608\,
            I => \il_min_comp2_D2\
        );

    \I__4511\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26599\
        );

    \I__4510\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26596\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__26599\,
            I => \N__26593\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__26596\,
            I => \N__26587\
        );

    \I__4507\ : Span4Mux_s2_v
    port map (
            O => \N__26593\,
            I => \N__26584\
        );

    \I__4506\ : CascadeMux
    port map (
            O => \N__26592\,
            I => \N__26581\
        );

    \I__4505\ : InMux
    port map (
            O => \N__26591\,
            I => \N__26577\
        );

    \I__4504\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26574\
        );

    \I__4503\ : Span4Mux_h
    port map (
            O => \N__26587\,
            I => \N__26569\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__26584\,
            I => \N__26569\
        );

    \I__4501\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26564\
        );

    \I__4500\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26564\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__26577\,
            I => \N__26559\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__26574\,
            I => \N__26559\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__26569\,
            I => \N__26556\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__26564\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__26559\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4494\ : Odrv4
    port map (
            O => \N__26556\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4493\ : IoInMux
    port map (
            O => \N__26549\,
            I => \N__26546\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__26546\,
            I => \N__26543\
        );

    \I__4491\ : Span4Mux_s2_v
    port map (
            O => \N__26543\,
            I => \N__26540\
        );

    \I__4490\ : Span4Mux_h
    port map (
            O => \N__26540\,
            I => \N__26537\
        );

    \I__4489\ : Span4Mux_v
    port map (
            O => \N__26537\,
            I => \N__26533\
        );

    \I__4488\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26530\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__26533\,
            I => \T23_c\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__26530\,
            I => \T23_c\
        );

    \I__4485\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26522\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__26522\,
            I => \N__26519\
        );

    \I__4483\ : Span4Mux_v
    port map (
            O => \N__26519\,
            I => \N__26516\
        );

    \I__4482\ : Span4Mux_v
    port map (
            O => \N__26516\,
            I => \N__26513\
        );

    \I__4481\ : Odrv4
    port map (
            O => \N__26513\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__4480\ : InMux
    port map (
            O => \N__26510\,
            I => \current_shift_inst.control_input_1_cry_3\
        );

    \I__4479\ : InMux
    port map (
            O => \N__26507\,
            I => \current_shift_inst.control_input_1_cry_4\
        );

    \I__4478\ : InMux
    port map (
            O => \N__26504\,
            I => \current_shift_inst.control_input_1_cry_5\
        );

    \I__4477\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26498\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__26498\,
            I => \N__26495\
        );

    \I__4475\ : Odrv12
    port map (
            O => \N__26495\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__4474\ : InMux
    port map (
            O => \N__26492\,
            I => \current_shift_inst.control_input_1_cry_6\
        );

    \I__4473\ : InMux
    port map (
            O => \N__26489\,
            I => \bfn_11_22_0_\
        );

    \I__4472\ : InMux
    port map (
            O => \N__26486\,
            I => \current_shift_inst.control_input_1_cry_8\
        );

    \I__4471\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26480\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__26480\,
            I => \N__26477\
        );

    \I__4469\ : Span12Mux_v
    port map (
            O => \N__26477\,
            I => \N__26474\
        );

    \I__4468\ : Odrv12
    port map (
            O => \N__26474\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__4467\ : InMux
    port map (
            O => \N__26471\,
            I => \current_shift_inst.control_input_1_cry_9\
        );

    \I__4466\ : InMux
    port map (
            O => \N__26468\,
            I => \current_shift_inst.control_input_1_cry_10\
        );

    \I__4465\ : InMux
    port map (
            O => \N__26465\,
            I => \N__26462\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__26462\,
            I => \current_shift_inst.control_input_1_axb_10\
        );

    \I__4463\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26456\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__26456\,
            I => \N__26453\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__26453\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__26450\,
            I => \phase_controller_inst2.start_timer_hc_RNOZ0Z_0_cascade_\
        );

    \I__4459\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26441\
        );

    \I__4458\ : InMux
    port map (
            O => \N__26446\,
            I => \N__26434\
        );

    \I__4457\ : InMux
    port map (
            O => \N__26445\,
            I => \N__26434\
        );

    \I__4456\ : InMux
    port map (
            O => \N__26444\,
            I => \N__26434\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__26441\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__26434\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__26429\,
            I => \phase_controller_inst2.start_timer_tr_0_sqmuxa_cascade_\
        );

    \I__4452\ : InMux
    port map (
            O => \N__26426\,
            I => \current_shift_inst.control_input_1_cry_0\
        );

    \I__4451\ : InMux
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__4449\ : Odrv12
    port map (
            O => \N__26417\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__4448\ : InMux
    port map (
            O => \N__26414\,
            I => \current_shift_inst.control_input_1_cry_1\
        );

    \I__4447\ : InMux
    port map (
            O => \N__26411\,
            I => \N__26408\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__26408\,
            I => \N__26405\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__26405\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__4444\ : InMux
    port map (
            O => \N__26402\,
            I => \current_shift_inst.control_input_1_cry_2\
        );

    \I__4443\ : InMux
    port map (
            O => \N__26399\,
            I => \N__26391\
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__26398\,
            I => \N__26386\
        );

    \I__4441\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26383\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__26396\,
            I => \N__26378\
        );

    \I__4439\ : CascadeMux
    port map (
            O => \N__26395\,
            I => \N__26375\
        );

    \I__4438\ : CascadeMux
    port map (
            O => \N__26394\,
            I => \N__26370\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__26391\,
            I => \N__26367\
        );

    \I__4436\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26364\
        );

    \I__4435\ : InMux
    port map (
            O => \N__26389\,
            I => \N__26361\
        );

    \I__4434\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26358\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__26383\,
            I => \N__26355\
        );

    \I__4432\ : CascadeMux
    port map (
            O => \N__26382\,
            I => \N__26352\
        );

    \I__4431\ : CascadeMux
    port map (
            O => \N__26381\,
            I => \N__26349\
        );

    \I__4430\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26345\
        );

    \I__4429\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26342\
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__26374\,
            I => \N__26335\
        );

    \I__4427\ : CascadeMux
    port map (
            O => \N__26373\,
            I => \N__26328\
        );

    \I__4426\ : InMux
    port map (
            O => \N__26370\,
            I => \N__26325\
        );

    \I__4425\ : Span4Mux_h
    port map (
            O => \N__26367\,
            I => \N__26322\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__26364\,
            I => \N__26317\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__26361\,
            I => \N__26317\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__26358\,
            I => \N__26314\
        );

    \I__4421\ : Span4Mux_h
    port map (
            O => \N__26355\,
            I => \N__26311\
        );

    \I__4420\ : InMux
    port map (
            O => \N__26352\,
            I => \N__26304\
        );

    \I__4419\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26304\
        );

    \I__4418\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26304\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__26345\,
            I => \N__26299\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__26342\,
            I => \N__26299\
        );

    \I__4415\ : InMux
    port map (
            O => \N__26341\,
            I => \N__26290\
        );

    \I__4414\ : InMux
    port map (
            O => \N__26340\,
            I => \N__26290\
        );

    \I__4413\ : InMux
    port map (
            O => \N__26339\,
            I => \N__26290\
        );

    \I__4412\ : InMux
    port map (
            O => \N__26338\,
            I => \N__26290\
        );

    \I__4411\ : InMux
    port map (
            O => \N__26335\,
            I => \N__26283\
        );

    \I__4410\ : InMux
    port map (
            O => \N__26334\,
            I => \N__26283\
        );

    \I__4409\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26283\
        );

    \I__4408\ : InMux
    port map (
            O => \N__26332\,
            I => \N__26276\
        );

    \I__4407\ : InMux
    port map (
            O => \N__26331\,
            I => \N__26276\
        );

    \I__4406\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26276\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__26325\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__26322\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__4403\ : Odrv12
    port map (
            O => \N__26317\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__4402\ : Odrv4
    port map (
            O => \N__26314\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__4401\ : Odrv4
    port map (
            O => \N__26311\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__26304\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__26299\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__26290\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__26283\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__26276\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__4395\ : CascadeMux
    port map (
            O => \N__26255\,
            I => \N__26252\
        );

    \I__4394\ : InMux
    port map (
            O => \N__26252\,
            I => \N__26249\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__26249\,
            I => \N__26245\
        );

    \I__4392\ : InMux
    port map (
            O => \N__26248\,
            I => \N__26241\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__26245\,
            I => \N__26238\
        );

    \I__4390\ : InMux
    port map (
            O => \N__26244\,
            I => \N__26235\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__26241\,
            I => \N__26232\
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__26238\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__26235\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__4386\ : Odrv4
    port map (
            O => \N__26232\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__4385\ : InMux
    port map (
            O => \N__26225\,
            I => \N__26221\
        );

    \I__4384\ : InMux
    port map (
            O => \N__26224\,
            I => \N__26218\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__26221\,
            I => \elapsed_time_ns_1_RNI81DJ11_0_2\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__26218\,
            I => \elapsed_time_ns_1_RNI81DJ11_0_2\
        );

    \I__4381\ : CascadeMux
    port map (
            O => \N__26213\,
            I => \elapsed_time_ns_1_RNI81DJ11_0_2_cascade_\
        );

    \I__4380\ : InMux
    port map (
            O => \N__26210\,
            I => \N__26206\
        );

    \I__4379\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26201\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__26206\,
            I => \N__26197\
        );

    \I__4377\ : InMux
    port map (
            O => \N__26205\,
            I => \N__26194\
        );

    \I__4376\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26191\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__26201\,
            I => \N__26188\
        );

    \I__4374\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26185\
        );

    \I__4373\ : Span4Mux_v
    port map (
            O => \N__26197\,
            I => \N__26180\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__26194\,
            I => \N__26180\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__26191\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3\
        );

    \I__4370\ : Odrv4
    port map (
            O => \N__26188\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__26185\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3\
        );

    \I__4368\ : Odrv4
    port map (
            O => \N__26180\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3\
        );

    \I__4367\ : InMux
    port map (
            O => \N__26171\,
            I => \N__26168\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__26168\,
            I => \phase_controller_inst1.stoper_hc.N_283\
        );

    \I__4365\ : CascadeMux
    port map (
            O => \N__26165\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_\
        );

    \I__4364\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26159\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__26159\,
            I => \N__26155\
        );

    \I__4362\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26152\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__26155\,
            I => \phase_controller_inst1.N_56\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__26152\,
            I => \phase_controller_inst1.N_56\
        );

    \I__4359\ : CascadeMux
    port map (
            O => \N__26147\,
            I => \N__26144\
        );

    \I__4358\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26138\
        );

    \I__4357\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26138\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__26138\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__4355\ : InMux
    port map (
            O => \N__26135\,
            I => \N__26132\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__26132\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__26129\,
            I => \N__26126\
        );

    \I__4352\ : InMux
    port map (
            O => \N__26126\,
            I => \N__26122\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__26125\,
            I => \N__26117\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__26122\,
            I => \N__26114\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__26121\,
            I => \N__26111\
        );

    \I__4348\ : InMux
    port map (
            O => \N__26120\,
            I => \N__26108\
        );

    \I__4347\ : InMux
    port map (
            O => \N__26117\,
            I => \N__26105\
        );

    \I__4346\ : Span4Mux_h
    port map (
            O => \N__26114\,
            I => \N__26102\
        );

    \I__4345\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26099\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__26108\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__26105\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4342\ : Odrv4
    port map (
            O => \N__26102\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__26099\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4340\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26087\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__26087\,
            I => \N__26084\
        );

    \I__4338\ : Span4Mux_h
    port map (
            O => \N__26084\,
            I => \N__26081\
        );

    \I__4337\ : Odrv4
    port map (
            O => \N__26081\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__26078\,
            I => \N__26073\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__26077\,
            I => \N__26069\
        );

    \I__4334\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26066\
        );

    \I__4333\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26063\
        );

    \I__4332\ : InMux
    port map (
            O => \N__26072\,
            I => \N__26058\
        );

    \I__4331\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26058\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__26066\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__26063\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__26058\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4327\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26048\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__26048\,
            I => \N__26045\
        );

    \I__4325\ : Span4Mux_v
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__26042\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__4323\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26026\
        );

    \I__4322\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26023\
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__26037\,
            I => \N__26019\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__26036\,
            I => \N__26016\
        );

    \I__4319\ : CascadeMux
    port map (
            O => \N__26035\,
            I => \N__26012\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__26034\,
            I => \N__26005\
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__26033\,
            I => \N__26000\
        );

    \I__4316\ : InMux
    port map (
            O => \N__26032\,
            I => \N__25987\
        );

    \I__4315\ : InMux
    port map (
            O => \N__26031\,
            I => \N__25987\
        );

    \I__4314\ : InMux
    port map (
            O => \N__26030\,
            I => \N__25987\
        );

    \I__4313\ : InMux
    port map (
            O => \N__26029\,
            I => \N__25987\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__26026\,
            I => \N__25982\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__26023\,
            I => \N__25982\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__26022\,
            I => \N__25978\
        );

    \I__4309\ : InMux
    port map (
            O => \N__26019\,
            I => \N__25961\
        );

    \I__4308\ : InMux
    port map (
            O => \N__26016\,
            I => \N__25961\
        );

    \I__4307\ : InMux
    port map (
            O => \N__26015\,
            I => \N__25961\
        );

    \I__4306\ : InMux
    port map (
            O => \N__26012\,
            I => \N__25961\
        );

    \I__4305\ : InMux
    port map (
            O => \N__26011\,
            I => \N__25961\
        );

    \I__4304\ : InMux
    port map (
            O => \N__26010\,
            I => \N__25961\
        );

    \I__4303\ : InMux
    port map (
            O => \N__26009\,
            I => \N__25961\
        );

    \I__4302\ : InMux
    port map (
            O => \N__26008\,
            I => \N__25961\
        );

    \I__4301\ : InMux
    port map (
            O => \N__26005\,
            I => \N__25944\
        );

    \I__4300\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25944\
        );

    \I__4299\ : InMux
    port map (
            O => \N__26003\,
            I => \N__25944\
        );

    \I__4298\ : InMux
    port map (
            O => \N__26000\,
            I => \N__25944\
        );

    \I__4297\ : InMux
    port map (
            O => \N__25999\,
            I => \N__25944\
        );

    \I__4296\ : InMux
    port map (
            O => \N__25998\,
            I => \N__25944\
        );

    \I__4295\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25944\
        );

    \I__4294\ : InMux
    port map (
            O => \N__25996\,
            I => \N__25944\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__25987\,
            I => \N__25941\
        );

    \I__4292\ : Span4Mux_v
    port map (
            O => \N__25982\,
            I => \N__25926\
        );

    \I__4291\ : InMux
    port map (
            O => \N__25981\,
            I => \N__25921\
        );

    \I__4290\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25921\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__25961\,
            I => \N__25918\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__25944\,
            I => \N__25915\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__25941\,
            I => \N__25912\
        );

    \I__4286\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25906\
        );

    \I__4285\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25906\
        );

    \I__4284\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25893\
        );

    \I__4283\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25893\
        );

    \I__4282\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25893\
        );

    \I__4281\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25893\
        );

    \I__4280\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25893\
        );

    \I__4279\ : InMux
    port map (
            O => \N__25933\,
            I => \N__25893\
        );

    \I__4278\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25884\
        );

    \I__4277\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25884\
        );

    \I__4276\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25884\
        );

    \I__4275\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25884\
        );

    \I__4274\ : Span4Mux_h
    port map (
            O => \N__25926\,
            I => \N__25881\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__25921\,
            I => \N__25876\
        );

    \I__4272\ : Span4Mux_v
    port map (
            O => \N__25918\,
            I => \N__25876\
        );

    \I__4271\ : Span4Mux_h
    port map (
            O => \N__25915\,
            I => \N__25873\
        );

    \I__4270\ : Span4Mux_h
    port map (
            O => \N__25912\,
            I => \N__25870\
        );

    \I__4269\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25867\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__25906\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__25893\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__25884\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4265\ : Odrv4
    port map (
            O => \N__25881\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4264\ : Odrv4
    port map (
            O => \N__25876\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4263\ : Odrv4
    port map (
            O => \N__25873\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__25870\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__25867\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4260\ : InMux
    port map (
            O => \N__25850\,
            I => \N__25847\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__25847\,
            I => \N__25842\
        );

    \I__4258\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25839\
        );

    \I__4257\ : InMux
    port map (
            O => \N__25845\,
            I => \N__25836\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__25842\,
            I => \elapsed_time_ns_1_RNIDP2KD1_0_1\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__25839\,
            I => \elapsed_time_ns_1_RNIDP2KD1_0_1\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__25836\,
            I => \elapsed_time_ns_1_RNIDP2KD1_0_1\
        );

    \I__4253\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25825\
        );

    \I__4252\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25822\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__25825\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_0_1Z0Z_1\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__25822\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_0_1Z0Z_1\
        );

    \I__4249\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25814\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__25814\,
            I => \N__25811\
        );

    \I__4247\ : Span4Mux_h
    port map (
            O => \N__25811\,
            I => \N__25808\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__25808\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__4245\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25801\
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__25804\,
            I => \N__25793\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__25801\,
            I => \N__25782\
        );

    \I__4242\ : InMux
    port map (
            O => \N__25800\,
            I => \N__25777\
        );

    \I__4241\ : InMux
    port map (
            O => \N__25799\,
            I => \N__25777\
        );

    \I__4240\ : InMux
    port map (
            O => \N__25798\,
            I => \N__25766\
        );

    \I__4239\ : InMux
    port map (
            O => \N__25797\,
            I => \N__25766\
        );

    \I__4238\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25766\
        );

    \I__4237\ : InMux
    port map (
            O => \N__25793\,
            I => \N__25766\
        );

    \I__4236\ : InMux
    port map (
            O => \N__25792\,
            I => \N__25766\
        );

    \I__4235\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25761\
        );

    \I__4234\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25761\
        );

    \I__4233\ : InMux
    port map (
            O => \N__25789\,
            I => \N__25752\
        );

    \I__4232\ : InMux
    port map (
            O => \N__25788\,
            I => \N__25752\
        );

    \I__4231\ : InMux
    port map (
            O => \N__25787\,
            I => \N__25752\
        );

    \I__4230\ : InMux
    port map (
            O => \N__25786\,
            I => \N__25752\
        );

    \I__4229\ : InMux
    port map (
            O => \N__25785\,
            I => \N__25749\
        );

    \I__4228\ : Span4Mux_h
    port map (
            O => \N__25782\,
            I => \N__25746\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__25777\,
            I => \phase_controller_inst1.stoper_hc.N_325\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__25766\,
            I => \phase_controller_inst1.stoper_hc.N_325\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__25761\,
            I => \phase_controller_inst1.stoper_hc.N_325\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__25752\,
            I => \phase_controller_inst1.stoper_hc.N_325\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__25749\,
            I => \phase_controller_inst1.stoper_hc.N_325\
        );

    \I__4222\ : Odrv4
    port map (
            O => \N__25746\,
            I => \phase_controller_inst1.stoper_hc.N_325\
        );

    \I__4221\ : CascadeMux
    port map (
            O => \N__25733\,
            I => \N__25725\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__25732\,
            I => \N__25722\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__25731\,
            I => \N__25716\
        );

    \I__4218\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25711\
        );

    \I__4217\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25706\
        );

    \I__4216\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25706\
        );

    \I__4215\ : InMux
    port map (
            O => \N__25725\,
            I => \N__25703\
        );

    \I__4214\ : InMux
    port map (
            O => \N__25722\,
            I => \N__25700\
        );

    \I__4213\ : InMux
    port map (
            O => \N__25721\,
            I => \N__25689\
        );

    \I__4212\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25689\
        );

    \I__4211\ : InMux
    port map (
            O => \N__25719\,
            I => \N__25689\
        );

    \I__4210\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25689\
        );

    \I__4209\ : InMux
    port map (
            O => \N__25715\,
            I => \N__25689\
        );

    \I__4208\ : InMux
    port map (
            O => \N__25714\,
            I => \N__25686\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__25711\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__25706\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__25703\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__25700\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__25689\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__25686\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__4201\ : InMux
    port map (
            O => \N__25673\,
            I => \N__25669\
        );

    \I__4200\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25666\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__25669\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_0_0Z0Z_3\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__25666\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_0_0Z0Z_3\
        );

    \I__4197\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25658\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__25658\,
            I => \N__25655\
        );

    \I__4195\ : Span4Mux_v
    port map (
            O => \N__25655\,
            I => \N__25652\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__25652\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__4193\ : CEMux
    port map (
            O => \N__25649\,
            I => \N__25646\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__25646\,
            I => \N__25643\
        );

    \I__4191\ : Span4Mux_v
    port map (
            O => \N__25643\,
            I => \N__25638\
        );

    \I__4190\ : CEMux
    port map (
            O => \N__25642\,
            I => \N__25635\
        );

    \I__4189\ : CEMux
    port map (
            O => \N__25641\,
            I => \N__25632\
        );

    \I__4188\ : Span4Mux_v
    port map (
            O => \N__25638\,
            I => \N__25629\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__25635\,
            I => \N__25626\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__25632\,
            I => \N__25623\
        );

    \I__4185\ : Span4Mux_h
    port map (
            O => \N__25629\,
            I => \N__25618\
        );

    \I__4184\ : Span4Mux_v
    port map (
            O => \N__25626\,
            I => \N__25618\
        );

    \I__4183\ : Span12Mux_s10_h
    port map (
            O => \N__25623\,
            I => \N__25615\
        );

    \I__4182\ : Span4Mux_h
    port map (
            O => \N__25618\,
            I => \N__25612\
        );

    \I__4181\ : Odrv12
    port map (
            O => \N__25615\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa_0\
        );

    \I__4180\ : Odrv4
    port map (
            O => \N__25612\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa_0\
        );

    \I__4179\ : CEMux
    port map (
            O => \N__25607\,
            I => \N__25603\
        );

    \I__4178\ : CEMux
    port map (
            O => \N__25606\,
            I => \N__25600\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__25603\,
            I => \N__25597\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__25600\,
            I => \N__25592\
        );

    \I__4175\ : Span4Mux_v
    port map (
            O => \N__25597\,
            I => \N__25589\
        );

    \I__4174\ : CEMux
    port map (
            O => \N__25596\,
            I => \N__25586\
        );

    \I__4173\ : CEMux
    port map (
            O => \N__25595\,
            I => \N__25583\
        );

    \I__4172\ : Span4Mux_v
    port map (
            O => \N__25592\,
            I => \N__25576\
        );

    \I__4171\ : Span4Mux_h
    port map (
            O => \N__25589\,
            I => \N__25576\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__25586\,
            I => \N__25576\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__25583\,
            I => \N__25573\
        );

    \I__4168\ : Span4Mux_h
    port map (
            O => \N__25576\,
            I => \N__25570\
        );

    \I__4167\ : Span4Mux_h
    port map (
            O => \N__25573\,
            I => \N__25567\
        );

    \I__4166\ : Odrv4
    port map (
            O => \N__25570\,
            I => \delay_measurement_inst.delay_hc_timer.N_433_i\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__25567\,
            I => \delay_measurement_inst.delay_hc_timer.N_433_i\
        );

    \I__4164\ : CascadeMux
    port map (
            O => \N__25562\,
            I => \N__25559\
        );

    \I__4163\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25556\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__25556\,
            I => \N__25553\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__25553\,
            I => \N__25550\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__25550\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__25547\,
            I => \N__25544\
        );

    \I__4158\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25541\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__25541\,
            I => \N__25538\
        );

    \I__4156\ : Span4Mux_h
    port map (
            O => \N__25538\,
            I => \N__25533\
        );

    \I__4155\ : InMux
    port map (
            O => \N__25537\,
            I => \N__25528\
        );

    \I__4154\ : InMux
    port map (
            O => \N__25536\,
            I => \N__25528\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__25533\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__25528\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__4151\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25520\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__25520\,
            I => \N__25516\
        );

    \I__4149\ : InMux
    port map (
            O => \N__25519\,
            I => \N__25512\
        );

    \I__4148\ : Span4Mux_h
    port map (
            O => \N__25516\,
            I => \N__25509\
        );

    \I__4147\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25506\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__25512\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7\
        );

    \I__4145\ : Odrv4
    port map (
            O => \N__25509\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__25506\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__25499\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7_cascade_\
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__25496\,
            I => \N__25493\
        );

    \I__4141\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25490\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__25490\,
            I => \N__25487\
        );

    \I__4139\ : Span4Mux_h
    port map (
            O => \N__25487\,
            I => \N__25483\
        );

    \I__4138\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25480\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__25483\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__25480\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__4135\ : CascadeMux
    port map (
            O => \N__25475\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\
        );

    \I__4134\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25469\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__25469\,
            I => \N__25465\
        );

    \I__4132\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25460\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__25465\,
            I => \N__25457\
        );

    \I__4130\ : InMux
    port map (
            O => \N__25464\,
            I => \N__25454\
        );

    \I__4129\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25451\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__25460\,
            I => \N__25445\
        );

    \I__4127\ : Span4Mux_h
    port map (
            O => \N__25457\,
            I => \N__25442\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__25454\,
            I => \N__25437\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__25451\,
            I => \N__25437\
        );

    \I__4124\ : InMux
    port map (
            O => \N__25450\,
            I => \N__25432\
        );

    \I__4123\ : InMux
    port map (
            O => \N__25449\,
            I => \N__25432\
        );

    \I__4122\ : InMux
    port map (
            O => \N__25448\,
            I => \N__25429\
        );

    \I__4121\ : Odrv4
    port map (
            O => \N__25445\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__4120\ : Odrv4
    port map (
            O => \N__25442\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__25437\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__25432\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__25429\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__4116\ : CascadeMux
    port map (
            O => \N__25418\,
            I => \elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_\
        );

    \I__4115\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25412\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__25412\,
            I => \N__25409\
        );

    \I__4113\ : Span4Mux_v
    port map (
            O => \N__25409\,
            I => \N__25406\
        );

    \I__4112\ : Odrv4
    port map (
            O => \N__25406\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__25403\,
            I => \N__25399\
        );

    \I__4110\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25396\
        );

    \I__4109\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25393\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__25396\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_0Z0Z_2\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__25393\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_0Z0Z_2\
        );

    \I__4106\ : InMux
    port map (
            O => \N__25388\,
            I => \N__25385\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__25385\,
            I => \N__25382\
        );

    \I__4104\ : Span4Mux_h
    port map (
            O => \N__25382\,
            I => \N__25379\
        );

    \I__4103\ : Odrv4
    port map (
            O => \N__25379\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__25376\,
            I => \N__25373\
        );

    \I__4101\ : InMux
    port map (
            O => \N__25373\,
            I => \N__25369\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__25372\,
            I => \N__25365\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__25369\,
            I => \N__25362\
        );

    \I__4098\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25358\
        );

    \I__4097\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25355\
        );

    \I__4096\ : Span4Mux_h
    port map (
            O => \N__25362\,
            I => \N__25352\
        );

    \I__4095\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25349\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__25358\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__25355\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__25352\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__25349\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4\
        );

    \I__4090\ : InMux
    port map (
            O => \N__25340\,
            I => \N__25337\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__25337\,
            I => \N__25334\
        );

    \I__4088\ : Span4Mux_h
    port map (
            O => \N__25334\,
            I => \N__25331\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__25331\,
            I => \N__25328\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__25328\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__4085\ : InMux
    port map (
            O => \N__25325\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__4084\ : InMux
    port map (
            O => \N__25322\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__4083\ : InMux
    port map (
            O => \N__25319\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__4082\ : InMux
    port map (
            O => \N__25316\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__4081\ : InMux
    port map (
            O => \N__25313\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__4080\ : InMux
    port map (
            O => \N__25310\,
            I => \bfn_11_15_0_\
        );

    \I__4079\ : InMux
    port map (
            O => \N__25307\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__4078\ : InMux
    port map (
            O => \N__25304\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__4077\ : InMux
    port map (
            O => \N__25301\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__4076\ : InMux
    port map (
            O => \N__25298\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__4075\ : InMux
    port map (
            O => \N__25295\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__4074\ : InMux
    port map (
            O => \N__25292\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__4073\ : InMux
    port map (
            O => \N__25289\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__4072\ : InMux
    port map (
            O => \N__25286\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__4071\ : InMux
    port map (
            O => \N__25283\,
            I => \bfn_11_14_0_\
        );

    \I__4070\ : InMux
    port map (
            O => \N__25280\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__4069\ : InMux
    port map (
            O => \N__25277\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__4068\ : InMux
    port map (
            O => \N__25274\,
            I => \N__25271\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__25271\,
            I => \N__25268\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__25268\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__4065\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25262\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__25262\,
            I => \N__25259\
        );

    \I__4063\ : Odrv12
    port map (
            O => \N__25259\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__4062\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25252\
        );

    \I__4061\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25249\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__25252\,
            I => \N__25245\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__25249\,
            I => \N__25241\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__25248\,
            I => \N__25236\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__25245\,
            I => \N__25231\
        );

    \I__4056\ : InMux
    port map (
            O => \N__25244\,
            I => \N__25228\
        );

    \I__4055\ : Span4Mux_v
    port map (
            O => \N__25241\,
            I => \N__25225\
        );

    \I__4054\ : InMux
    port map (
            O => \N__25240\,
            I => \N__25214\
        );

    \I__4053\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25214\
        );

    \I__4052\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25214\
        );

    \I__4051\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25214\
        );

    \I__4050\ : InMux
    port map (
            O => \N__25234\,
            I => \N__25214\
        );

    \I__4049\ : Span4Mux_v
    port map (
            O => \N__25231\,
            I => \N__25211\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__25228\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__25225\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__25214\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__25211\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__4044\ : InMux
    port map (
            O => \N__25202\,
            I => \N__25196\
        );

    \I__4043\ : InMux
    port map (
            O => \N__25201\,
            I => \N__25191\
        );

    \I__4042\ : InMux
    port map (
            O => \N__25200\,
            I => \N__25188\
        );

    \I__4041\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25185\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__25196\,
            I => \N__25182\
        );

    \I__4039\ : InMux
    port map (
            O => \N__25195\,
            I => \N__25177\
        );

    \I__4038\ : InMux
    port map (
            O => \N__25194\,
            I => \N__25177\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__25191\,
            I => \N__25174\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__25188\,
            I => \N__25171\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__25185\,
            I => \N__25164\
        );

    \I__4034\ : Span4Mux_h
    port map (
            O => \N__25182\,
            I => \N__25164\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25164\
        );

    \I__4032\ : Odrv4
    port map (
            O => \N__25174\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__4031\ : Odrv12
    port map (
            O => \N__25171\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__4030\ : Odrv4
    port map (
            O => \N__25164\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__25157\,
            I => \N__25154\
        );

    \I__4028\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25151\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__25151\,
            I => \N__25147\
        );

    \I__4026\ : InMux
    port map (
            O => \N__25150\,
            I => \N__25143\
        );

    \I__4025\ : Span4Mux_h
    port map (
            O => \N__25147\,
            I => \N__25140\
        );

    \I__4024\ : InMux
    port map (
            O => \N__25146\,
            I => \N__25137\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__25143\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__25140\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__25137\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4020\ : SRMux
    port map (
            O => \N__25130\,
            I => \N__25127\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__25127\,
            I => \N__25122\
        );

    \I__4018\ : SRMux
    port map (
            O => \N__25126\,
            I => \N__25119\
        );

    \I__4017\ : SRMux
    port map (
            O => \N__25125\,
            I => \N__25115\
        );

    \I__4016\ : Span4Mux_h
    port map (
            O => \N__25122\,
            I => \N__25110\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__25119\,
            I => \N__25110\
        );

    \I__4014\ : SRMux
    port map (
            O => \N__25118\,
            I => \N__25107\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__25115\,
            I => \N__25104\
        );

    \I__4012\ : Span4Mux_v
    port map (
            O => \N__25110\,
            I => \N__25101\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__25107\,
            I => \N__25098\
        );

    \I__4010\ : Span4Mux_h
    port map (
            O => \N__25104\,
            I => \N__25095\
        );

    \I__4009\ : Span4Mux_h
    port map (
            O => \N__25101\,
            I => \N__25090\
        );

    \I__4008\ : Span4Mux_v
    port map (
            O => \N__25098\,
            I => \N__25090\
        );

    \I__4007\ : Sp12to4
    port map (
            O => \N__25095\,
            I => \N__25087\
        );

    \I__4006\ : Span4Mux_h
    port map (
            O => \N__25090\,
            I => \N__25084\
        );

    \I__4005\ : Odrv12
    port map (
            O => \N__25087\,
            I => \phase_controller_inst1.stoper_hc.un1_stoper_state12_1_0_i\
        );

    \I__4004\ : Odrv4
    port map (
            O => \N__25084\,
            I => \phase_controller_inst1.stoper_hc.un1_stoper_state12_1_0_i\
        );

    \I__4003\ : InMux
    port map (
            O => \N__25079\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__4002\ : IoInMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__4000\ : Span4Mux_s3_v
    port map (
            O => \N__25070\,
            I => \N__25067\
        );

    \I__3999\ : Sp12to4
    port map (
            O => \N__25067\,
            I => \N__25064\
        );

    \I__3998\ : Span12Mux_h
    port map (
            O => \N__25064\,
            I => \N__25060\
        );

    \I__3997\ : InMux
    port map (
            O => \N__25063\,
            I => \N__25057\
        );

    \I__3996\ : Odrv12
    port map (
            O => \N__25060\,
            I => \T12_c\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__25057\,
            I => \T12_c\
        );

    \I__3994\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25046\
        );

    \I__3993\ : InMux
    port map (
            O => \N__25051\,
            I => \N__25046\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__25046\,
            I => state_ns_i_a3_1
        );

    \I__3991\ : ClkMux
    port map (
            O => \N__25043\,
            I => \N__25037\
        );

    \I__3990\ : ClkMux
    port map (
            O => \N__25042\,
            I => \N__25037\
        );

    \I__3989\ : GlobalMux
    port map (
            O => \N__25037\,
            I => \N__25034\
        );

    \I__3988\ : gio2CtrlBuf
    port map (
            O => \N__25034\,
            I => delay_hc_input_c_g
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__25031\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__3986\ : InMux
    port map (
            O => \N__25028\,
            I => \N__25025\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__25025\,
            I => \N__25022\
        );

    \I__3984\ : Span4Mux_v
    port map (
            O => \N__25022\,
            I => \N__25019\
        );

    \I__3983\ : Odrv4
    port map (
            O => \N__25019\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__25016\,
            I => \N__25013\
        );

    \I__3981\ : InMux
    port map (
            O => \N__25013\,
            I => \N__25010\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__25010\,
            I => \N__25007\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__25007\,
            I => \N__25004\
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__25004\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0\
        );

    \I__3977\ : CascadeMux
    port map (
            O => \N__25001\,
            I => \phase_controller_inst1.stoper_hc.N_45_cascade_\
        );

    \I__3976\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24991\
        );

    \I__3975\ : InMux
    port map (
            O => \N__24997\,
            I => \N__24982\
        );

    \I__3974\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24982\
        );

    \I__3973\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24982\
        );

    \I__3972\ : InMux
    port map (
            O => \N__24994\,
            I => \N__24982\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__24991\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__24982\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3969\ : CascadeMux
    port map (
            O => \N__24977\,
            I => \N__24972\
        );

    \I__3968\ : CascadeMux
    port map (
            O => \N__24976\,
            I => \N__24966\
        );

    \I__3967\ : CascadeMux
    port map (
            O => \N__24975\,
            I => \N__24963\
        );

    \I__3966\ : InMux
    port map (
            O => \N__24972\,
            I => \N__24954\
        );

    \I__3965\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24954\
        );

    \I__3964\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24954\
        );

    \I__3963\ : InMux
    port map (
            O => \N__24969\,
            I => \N__24954\
        );

    \I__3962\ : InMux
    port map (
            O => \N__24966\,
            I => \N__24951\
        );

    \I__3961\ : InMux
    port map (
            O => \N__24963\,
            I => \N__24948\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__24954\,
            I => \N__24945\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__24951\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__24948\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__24945\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__24938\,
            I => \N__24934\
        );

    \I__3955\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24931\
        );

    \I__3954\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24928\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__24931\,
            I => \N__24922\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__24928\,
            I => \N__24922\
        );

    \I__3951\ : InMux
    port map (
            O => \N__24927\,
            I => \N__24919\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__24922\,
            I => \N__24914\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__24919\,
            I => \N__24914\
        );

    \I__3948\ : Span4Mux_h
    port map (
            O => \N__24914\,
            I => \N__24911\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__24911\,
            I => \il_max_comp2_D2\
        );

    \I__3946\ : CascadeMux
    port map (
            O => \N__24908\,
            I => \phase_controller_inst1.stoper_hc.N_325_cascade_\
        );

    \I__3945\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24902\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__24902\,
            I => \N__24899\
        );

    \I__3943\ : Span4Mux_h
    port map (
            O => \N__24899\,
            I => \N__24896\
        );

    \I__3942\ : Odrv4
    port map (
            O => \N__24896\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__24893\,
            I => \N__24888\
        );

    \I__3940\ : InMux
    port map (
            O => \N__24892\,
            I => \N__24884\
        );

    \I__3939\ : InMux
    port map (
            O => \N__24891\,
            I => \N__24878\
        );

    \I__3938\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24875\
        );

    \I__3937\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24872\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__24884\,
            I => \N__24869\
        );

    \I__3935\ : InMux
    port map (
            O => \N__24883\,
            I => \N__24865\
        );

    \I__3934\ : InMux
    port map (
            O => \N__24882\,
            I => \N__24861\
        );

    \I__3933\ : InMux
    port map (
            O => \N__24881\,
            I => \N__24858\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__24878\,
            I => \N__24855\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__24875\,
            I => \N__24850\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__24872\,
            I => \N__24850\
        );

    \I__3929\ : Span4Mux_v
    port map (
            O => \N__24869\,
            I => \N__24847\
        );

    \I__3928\ : InMux
    port map (
            O => \N__24868\,
            I => \N__24844\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__24865\,
            I => \N__24841\
        );

    \I__3926\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24838\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__24861\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__24858\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__3923\ : Odrv4
    port map (
            O => \N__24855\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__24850\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__24847\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__24844\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__24841\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__24838\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__24821\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2_cascade_\
        );

    \I__3916\ : CascadeMux
    port map (
            O => \N__24818\,
            I => \phase_controller_inst1.stoper_hc.N_307_cascade_\
        );

    \I__3915\ : CascadeMux
    port map (
            O => \N__24815\,
            I => \N__24812\
        );

    \I__3914\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24806\
        );

    \I__3912\ : Span4Mux_h
    port map (
            O => \N__24806\,
            I => \N__24801\
        );

    \I__3911\ : InMux
    port map (
            O => \N__24805\,
            I => \N__24796\
        );

    \I__3910\ : InMux
    port map (
            O => \N__24804\,
            I => \N__24796\
        );

    \I__3909\ : Odrv4
    port map (
            O => \N__24801\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__24796\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__3907\ : CascadeMux
    port map (
            O => \N__24791\,
            I => \N__24788\
        );

    \I__3906\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24783\
        );

    \I__3905\ : InMux
    port map (
            O => \N__24787\,
            I => \N__24778\
        );

    \I__3904\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24778\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__24783\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__24778\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__24773\,
            I => \N__24768\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__24772\,
            I => \N__24765\
        );

    \I__3899\ : InMux
    port map (
            O => \N__24771\,
            I => \N__24762\
        );

    \I__3898\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24757\
        );

    \I__3897\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24757\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__24762\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1Z0Z_2\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__24757\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1Z0Z_2\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__24752\,
            I => \N__24745\
        );

    \I__3893\ : InMux
    port map (
            O => \N__24751\,
            I => \N__24728\
        );

    \I__3892\ : InMux
    port map (
            O => \N__24750\,
            I => \N__24728\
        );

    \I__3891\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24728\
        );

    \I__3890\ : InMux
    port map (
            O => \N__24748\,
            I => \N__24728\
        );

    \I__3889\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24715\
        );

    \I__3888\ : InMux
    port map (
            O => \N__24744\,
            I => \N__24715\
        );

    \I__3887\ : InMux
    port map (
            O => \N__24743\,
            I => \N__24715\
        );

    \I__3886\ : InMux
    port map (
            O => \N__24742\,
            I => \N__24715\
        );

    \I__3885\ : InMux
    port map (
            O => \N__24741\,
            I => \N__24715\
        );

    \I__3884\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24710\
        );

    \I__3883\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24710\
        );

    \I__3882\ : InMux
    port map (
            O => \N__24738\,
            I => \N__24705\
        );

    \I__3881\ : InMux
    port map (
            O => \N__24737\,
            I => \N__24705\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__24728\,
            I => \N__24702\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__24727\,
            I => \N__24696\
        );

    \I__3878\ : CascadeMux
    port map (
            O => \N__24726\,
            I => \N__24693\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__24715\,
            I => \N__24681\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__24710\,
            I => \N__24681\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__24705\,
            I => \N__24681\
        );

    \I__3874\ : Span4Mux_v
    port map (
            O => \N__24702\,
            I => \N__24678\
        );

    \I__3873\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24675\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__24700\,
            I => \N__24671\
        );

    \I__3871\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24651\
        );

    \I__3870\ : InMux
    port map (
            O => \N__24696\,
            I => \N__24651\
        );

    \I__3869\ : InMux
    port map (
            O => \N__24693\,
            I => \N__24651\
        );

    \I__3868\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24651\
        );

    \I__3867\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24651\
        );

    \I__3866\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24651\
        );

    \I__3865\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24651\
        );

    \I__3864\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24651\
        );

    \I__3863\ : Span4Mux_v
    port map (
            O => \N__24681\,
            I => \N__24646\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__24678\,
            I => \N__24646\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__24675\,
            I => \N__24643\
        );

    \I__3860\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24638\
        );

    \I__3859\ : InMux
    port map (
            O => \N__24671\,
            I => \N__24638\
        );

    \I__3858\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24631\
        );

    \I__3857\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24631\
        );

    \I__3856\ : InMux
    port map (
            O => \N__24668\,
            I => \N__24631\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__24651\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15\
        );

    \I__3854\ : Odrv4
    port map (
            O => \N__24646\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__24643\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__24638\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__24631\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15\
        );

    \I__3850\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__24617\,
            I => \N__24614\
        );

    \I__3848\ : Span4Mux_v
    port map (
            O => \N__24614\,
            I => \N__24611\
        );

    \I__3847\ : Span4Mux_h
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__24608\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__3845\ : InMux
    port map (
            O => \N__24605\,
            I => \N__24601\
        );

    \I__3844\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24598\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__24601\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__24598\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__24593\,
            I => \N__24590\
        );

    \I__3840\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24587\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__24587\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__3838\ : InMux
    port map (
            O => \N__24584\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__3837\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24578\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__24578\,
            I => \N__24575\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__24575\,
            I => \il_max_comp1_D1\
        );

    \I__3834\ : InMux
    port map (
            O => \N__24572\,
            I => \N__24568\
        );

    \I__3833\ : InMux
    port map (
            O => \N__24571\,
            I => \N__24565\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__24568\,
            I => \N__24561\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__24565\,
            I => \N__24558\
        );

    \I__3830\ : InMux
    port map (
            O => \N__24564\,
            I => \N__24555\
        );

    \I__3829\ : Span12Mux_h
    port map (
            O => \N__24561\,
            I => \N__24552\
        );

    \I__3828\ : Span4Mux_h
    port map (
            O => \N__24558\,
            I => \N__24547\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__24555\,
            I => \N__24547\
        );

    \I__3826\ : Odrv12
    port map (
            O => \N__24552\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__24547\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__3824\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__3822\ : Span4Mux_v
    port map (
            O => \N__24536\,
            I => \N__24533\
        );

    \I__3821\ : Odrv4
    port map (
            O => \N__24533\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\
        );

    \I__3820\ : InMux
    port map (
            O => \N__24530\,
            I => \N__24527\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__24527\,
            I => \N__24519\
        );

    \I__3818\ : InMux
    port map (
            O => \N__24526\,
            I => \N__24516\
        );

    \I__3817\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24511\
        );

    \I__3816\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24511\
        );

    \I__3815\ : InMux
    port map (
            O => \N__24523\,
            I => \N__24506\
        );

    \I__3814\ : InMux
    port map (
            O => \N__24522\,
            I => \N__24506\
        );

    \I__3813\ : Span4Mux_h
    port map (
            O => \N__24519\,
            I => \N__24503\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__24516\,
            I => \N__24500\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__24511\,
            I => \N__24495\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__24506\,
            I => \N__24495\
        );

    \I__3809\ : Span4Mux_v
    port map (
            O => \N__24503\,
            I => \N__24492\
        );

    \I__3808\ : Span4Mux_v
    port map (
            O => \N__24500\,
            I => \N__24487\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__24495\,
            I => \N__24487\
        );

    \I__3806\ : Odrv4
    port map (
            O => \N__24492\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__3805\ : Odrv4
    port map (
            O => \N__24487\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__3804\ : InMux
    port map (
            O => \N__24482\,
            I => \N__24475\
        );

    \I__3803\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24475\
        );

    \I__3802\ : InMux
    port map (
            O => \N__24480\,
            I => \N__24471\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__24475\,
            I => \N__24468\
        );

    \I__3800\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24465\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__24471\,
            I => \N__24461\
        );

    \I__3798\ : Span4Mux_h
    port map (
            O => \N__24468\,
            I => \N__24458\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__24465\,
            I => \N__24455\
        );

    \I__3796\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24452\
        );

    \I__3795\ : Odrv12
    port map (
            O => \N__24461\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19\
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__24458\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__24455\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__24452\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19\
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__24443\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_\
        );

    \I__3790\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24435\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__24439\,
            I => \N__24432\
        );

    \I__3788\ : InMux
    port map (
            O => \N__24438\,
            I => \N__24429\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__24435\,
            I => \N__24426\
        );

    \I__3786\ : InMux
    port map (
            O => \N__24432\,
            I => \N__24423\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__24429\,
            I => \N__24418\
        );

    \I__3784\ : Span4Mux_h
    port map (
            O => \N__24426\,
            I => \N__24418\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__24423\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a5_1_1_9\
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__24418\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a5_1_1_9\
        );

    \I__3781\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24410\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__24410\,
            I => \N__24405\
        );

    \I__3779\ : InMux
    port map (
            O => \N__24409\,
            I => \N__24401\
        );

    \I__3778\ : InMux
    port map (
            O => \N__24408\,
            I => \N__24398\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__24405\,
            I => \N__24395\
        );

    \I__3776\ : InMux
    port map (
            O => \N__24404\,
            I => \N__24392\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__24401\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__24398\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9\
        );

    \I__3773\ : Odrv4
    port map (
            O => \N__24395\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__24392\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9\
        );

    \I__3771\ : InMux
    port map (
            O => \N__24383\,
            I => \N__24380\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__24380\,
            I => \N__24377\
        );

    \I__3769\ : Odrv12
    port map (
            O => \N__24377\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1Z0Z_6\
        );

    \I__3768\ : InMux
    port map (
            O => \N__24374\,
            I => \N__24370\
        );

    \I__3767\ : InMux
    port map (
            O => \N__24373\,
            I => \N__24367\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__24370\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__24367\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3764\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24359\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24356\
        );

    \I__3762\ : Span4Mux_v
    port map (
            O => \N__24356\,
            I => \N__24353\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__24353\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__3760\ : CascadeMux
    port map (
            O => \N__24350\,
            I => \N__24347\
        );

    \I__3759\ : InMux
    port map (
            O => \N__24347\,
            I => \N__24344\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__24344\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__3757\ : InMux
    port map (
            O => \N__24341\,
            I => \N__24338\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__24338\,
            I => \N__24335\
        );

    \I__3755\ : Span4Mux_v
    port map (
            O => \N__24335\,
            I => \N__24332\
        );

    \I__3754\ : Sp12to4
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__3753\ : Odrv12
    port map (
            O => \N__24329\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__3752\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24322\
        );

    \I__3751\ : InMux
    port map (
            O => \N__24325\,
            I => \N__24319\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__24322\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__24319\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__3747\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24308\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__24308\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__3745\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24301\
        );

    \I__3744\ : InMux
    port map (
            O => \N__24304\,
            I => \N__24298\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__24301\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__24298\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__24293\,
            I => \N__24290\
        );

    \I__3740\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__24287\,
            I => \N__24284\
        );

    \I__3738\ : Odrv12
    port map (
            O => \N__24284\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__3737\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24278\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__24278\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__3735\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24272\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__24272\,
            I => \N__24269\
        );

    \I__3733\ : Span4Mux_h
    port map (
            O => \N__24269\,
            I => \N__24266\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__24266\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__3731\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24259\
        );

    \I__3730\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24256\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__24259\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__24256\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__3726\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24245\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__24245\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__3724\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24239\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__24239\,
            I => \N__24236\
        );

    \I__3722\ : Span4Mux_h
    port map (
            O => \N__24236\,
            I => \N__24233\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__24233\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__3720\ : InMux
    port map (
            O => \N__24230\,
            I => \N__24226\
        );

    \I__3719\ : InMux
    port map (
            O => \N__24229\,
            I => \N__24223\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__24226\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__24223\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__24218\,
            I => \N__24215\
        );

    \I__3715\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24212\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__24212\,
            I => \N__24209\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__24209\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__3712\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__24203\,
            I => \N__24200\
        );

    \I__3710\ : Span4Mux_h
    port map (
            O => \N__24200\,
            I => \N__24197\
        );

    \I__3709\ : Span4Mux_h
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__24194\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__3707\ : InMux
    port map (
            O => \N__24191\,
            I => \N__24187\
        );

    \I__3706\ : InMux
    port map (
            O => \N__24190\,
            I => \N__24184\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__24187\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__24184\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__24179\,
            I => \N__24176\
        );

    \I__3702\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24173\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__24173\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__3700\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24167\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__24167\,
            I => \N__24164\
        );

    \I__3698\ : Span4Mux_h
    port map (
            O => \N__24164\,
            I => \N__24161\
        );

    \I__3697\ : Span4Mux_h
    port map (
            O => \N__24161\,
            I => \N__24158\
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__24158\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__3695\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24151\
        );

    \I__3694\ : InMux
    port map (
            O => \N__24154\,
            I => \N__24148\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__24151\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__24148\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__24143\,
            I => \N__24140\
        );

    \I__3690\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24137\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__24137\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__3688\ : InMux
    port map (
            O => \N__24134\,
            I => \N__24130\
        );

    \I__3687\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24127\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__24130\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__24127\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__24122\,
            I => \N__24119\
        );

    \I__3683\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24116\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__24116\,
            I => \N__24113\
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__24113\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__3680\ : InMux
    port map (
            O => \N__24110\,
            I => \N__24106\
        );

    \I__3679\ : InMux
    port map (
            O => \N__24109\,
            I => \N__24103\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__24106\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__24103\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__24098\,
            I => \N__24095\
        );

    \I__3675\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24092\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__24092\,
            I => \N__24089\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__24089\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__3672\ : InMux
    port map (
            O => \N__24086\,
            I => \N__24082\
        );

    \I__3671\ : InMux
    port map (
            O => \N__24085\,
            I => \N__24079\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__24082\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__24079\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3668\ : CascadeMux
    port map (
            O => \N__24074\,
            I => \N__24071\
        );

    \I__3667\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24068\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__24068\,
            I => \N__24065\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__24065\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__3664\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24059\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__24059\,
            I => \N__24056\
        );

    \I__3662\ : Span4Mux_h
    port map (
            O => \N__24056\,
            I => \N__24053\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__24053\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__3660\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24046\
        );

    \I__3659\ : InMux
    port map (
            O => \N__24049\,
            I => \N__24043\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__24046\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__24043\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3656\ : CascadeMux
    port map (
            O => \N__24038\,
            I => \N__24035\
        );

    \I__3655\ : InMux
    port map (
            O => \N__24035\,
            I => \N__24032\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__24032\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__3653\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24025\
        );

    \I__3652\ : InMux
    port map (
            O => \N__24028\,
            I => \N__24022\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__24025\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__24022\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3649\ : CascadeMux
    port map (
            O => \N__24017\,
            I => \N__24014\
        );

    \I__3648\ : InMux
    port map (
            O => \N__24014\,
            I => \N__24011\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__24008\
        );

    \I__3646\ : Odrv4
    port map (
            O => \N__24008\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__3645\ : InMux
    port map (
            O => \N__24005\,
            I => \N__24002\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__24002\,
            I => \N__23999\
        );

    \I__3643\ : Span4Mux_v
    port map (
            O => \N__23999\,
            I => \N__23996\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__23996\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__3641\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23989\
        );

    \I__3640\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23986\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__23989\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__23986\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3637\ : CascadeMux
    port map (
            O => \N__23981\,
            I => \N__23978\
        );

    \I__3636\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23975\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__23975\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__3634\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23969\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__23969\,
            I => \N__23966\
        );

    \I__3632\ : Span4Mux_h
    port map (
            O => \N__23966\,
            I => \N__23963\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__23963\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__3630\ : InMux
    port map (
            O => \N__23960\,
            I => \N__23956\
        );

    \I__3629\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23953\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__23956\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__23953\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3626\ : CascadeMux
    port map (
            O => \N__23948\,
            I => \N__23945\
        );

    \I__3625\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23942\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__23942\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__3623\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23935\
        );

    \I__3622\ : InMux
    port map (
            O => \N__23938\,
            I => \N__23932\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__23935\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__23932\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3619\ : InMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__23924\,
            I => \N__23921\
        );

    \I__3617\ : Span4Mux_v
    port map (
            O => \N__23921\,
            I => \N__23918\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__23918\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__23915\,
            I => \N__23912\
        );

    \I__3614\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23909\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__23909\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__3612\ : IoInMux
    port map (
            O => \N__23906\,
            I => \N__23903\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__23903\,
            I => \N__23900\
        );

    \I__3610\ : Odrv4
    port map (
            O => \N__23900\,
            I => s3_phy_c
        );

    \I__3609\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23894\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__23894\,
            I => \N__23891\
        );

    \I__3607\ : Span4Mux_h
    port map (
            O => \N__23891\,
            I => \N__23888\
        );

    \I__3606\ : Span4Mux_v
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__3605\ : Odrv4
    port map (
            O => \N__23885\,
            I => il_min_comp1_c
        );

    \I__3604\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23876\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__23876\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__3601\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23870\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__23870\,
            I => \N__23867\
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__23867\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__3598\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23861\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__23861\,
            I => \N__23858\
        );

    \I__3596\ : Odrv12
    port map (
            O => \N__23858\,
            I => \il_min_comp1_D1\
        );

    \I__3595\ : InMux
    port map (
            O => \N__23855\,
            I => \N__23852\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__23852\,
            I => \N__23849\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__23849\,
            I => \N__23846\
        );

    \I__3592\ : Span4Mux_v
    port map (
            O => \N__23846\,
            I => \N__23843\
        );

    \I__3591\ : Span4Mux_v
    port map (
            O => \N__23843\,
            I => \N__23840\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__23840\,
            I => il_max_comp1_c
        );

    \I__3589\ : CascadeMux
    port map (
            O => \N__23837\,
            I => \N__23834\
        );

    \I__3588\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23831\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__23831\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__3586\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23824\
        );

    \I__3585\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23821\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__23824\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__23821\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__23816\,
            I => \N__23813\
        );

    \I__3581\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23810\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__23810\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__3579\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23803\
        );

    \I__3578\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23800\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__23803\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__23800\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__23795\,
            I => \N__23792\
        );

    \I__3574\ : InMux
    port map (
            O => \N__23792\,
            I => \N__23789\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__23789\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__3572\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23782\
        );

    \I__3571\ : InMux
    port map (
            O => \N__23785\,
            I => \N__23779\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__23782\,
            I => \N__23776\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__23779\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__23776\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4\
        );

    \I__3567\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23768\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__23768\,
            I => \N__23763\
        );

    \I__3565\ : InMux
    port map (
            O => \N__23767\,
            I => \N__23758\
        );

    \I__3564\ : InMux
    port map (
            O => \N__23766\,
            I => \N__23758\
        );

    \I__3563\ : Odrv4
    port map (
            O => \N__23763\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__23758\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\
        );

    \I__3561\ : InMux
    port map (
            O => \N__23753\,
            I => \N__23749\
        );

    \I__3560\ : InMux
    port map (
            O => \N__23752\,
            I => \N__23746\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__23749\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__23746\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\
        );

    \I__3557\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23736\
        );

    \I__3556\ : InMux
    port map (
            O => \N__23740\,
            I => \N__23731\
        );

    \I__3555\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23731\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__23736\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__23731\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__23726\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__23723\,
            I => \N__23719\
        );

    \I__3550\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23716\
        );

    \I__3549\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23713\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__23716\,
            I => \N__23707\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__23713\,
            I => \N__23707\
        );

    \I__3546\ : InMux
    port map (
            O => \N__23712\,
            I => \N__23704\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__23707\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__23704\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__23699\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__23696\,
            I => \N__23692\
        );

    \I__3541\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23688\
        );

    \I__3540\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23685\
        );

    \I__3539\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23682\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__23688\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__23685\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__23682\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__23675\,
            I => \N__23671\
        );

    \I__3534\ : InMux
    port map (
            O => \N__23674\,
            I => \N__23667\
        );

    \I__3533\ : InMux
    port map (
            O => \N__23671\,
            I => \N__23664\
        );

    \I__3532\ : InMux
    port map (
            O => \N__23670\,
            I => \N__23661\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__23667\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__23664\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__23661\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__3528\ : CEMux
    port map (
            O => \N__23654\,
            I => \N__23639\
        );

    \I__3527\ : CEMux
    port map (
            O => \N__23653\,
            I => \N__23639\
        );

    \I__3526\ : CEMux
    port map (
            O => \N__23652\,
            I => \N__23639\
        );

    \I__3525\ : CEMux
    port map (
            O => \N__23651\,
            I => \N__23639\
        );

    \I__3524\ : CEMux
    port map (
            O => \N__23650\,
            I => \N__23639\
        );

    \I__3523\ : GlobalMux
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__3522\ : gio2CtrlBuf
    port map (
            O => \N__23636\,
            I => \delay_measurement_inst.delay_hc_timer.N_432_i_g\
        );

    \I__3521\ : IoInMux
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__3519\ : Span4Mux_s0_v
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__3518\ : Span4Mux_h
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__3517\ : Span4Mux_v
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__3516\ : Span4Mux_v
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__3515\ : Odrv4
    port map (
            O => \N__23615\,
            I => \delay_measurement_inst.delay_hc_timer.N_432_i\
        );

    \I__3514\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__23609\,
            I => \N__23606\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__23606\,
            I => \N__23603\
        );

    \I__3511\ : Span4Mux_v
    port map (
            O => \N__23603\,
            I => \N__23600\
        );

    \I__3510\ : Span4Mux_v
    port map (
            O => \N__23600\,
            I => \N__23597\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__23597\,
            I => \il_min_comp2_D1\
        );

    \I__3508\ : InMux
    port map (
            O => \N__23594\,
            I => \N__23591\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__23591\,
            I => \N__23587\
        );

    \I__3506\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23584\
        );

    \I__3505\ : Span4Mux_h
    port map (
            O => \N__23587\,
            I => \N__23581\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__23584\,
            I => \N__23578\
        );

    \I__3503\ : Odrv4
    port map (
            O => \N__23581\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__3502\ : Odrv12
    port map (
            O => \N__23578\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__3500\ : InMux
    port map (
            O => \N__23570\,
            I => \N__23567\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__23567\,
            I => \elapsed_time_ns_1_RNIT6ND11_0_25\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__23564\,
            I => \elapsed_time_ns_1_RNIT6ND11_0_25_cascade_\
        );

    \I__3497\ : InMux
    port map (
            O => \N__23561\,
            I => \N__23558\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__23558\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_o5_6Z0Z_15\
        );

    \I__3495\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23551\
        );

    \I__3494\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23548\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__23551\,
            I => \N__23543\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__23548\,
            I => \N__23543\
        );

    \I__3491\ : Span4Mux_h
    port map (
            O => \N__23543\,
            I => \N__23540\
        );

    \I__3490\ : Odrv4
    port map (
            O => \N__23540\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__3489\ : InMux
    port map (
            O => \N__23537\,
            I => \N__23531\
        );

    \I__3488\ : InMux
    port map (
            O => \N__23536\,
            I => \N__23531\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__23531\,
            I => \elapsed_time_ns_1_RNIV8ND11_0_27\
        );

    \I__3486\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23524\
        );

    \I__3485\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23521\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__23524\,
            I => \N__23516\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__23521\,
            I => \N__23516\
        );

    \I__3482\ : Span4Mux_h
    port map (
            O => \N__23516\,
            I => \N__23513\
        );

    \I__3481\ : Odrv4
    port map (
            O => \N__23513\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__3480\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23504\
        );

    \I__3479\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23504\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__23504\,
            I => \elapsed_time_ns_1_RNIU7ND11_0_26\
        );

    \I__3477\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23498\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__23498\,
            I => \N__23494\
        );

    \I__3475\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23491\
        );

    \I__3474\ : Span4Mux_h
    port map (
            O => \N__23494\,
            I => \N__23488\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__23491\,
            I => \N__23485\
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__23488\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__3471\ : Odrv12
    port map (
            O => \N__23485\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__23480\,
            I => \N__23477\
        );

    \I__3469\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23473\
        );

    \I__3468\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23470\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__23473\,
            I => \elapsed_time_ns_1_RNI0AND11_0_28\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__23470\,
            I => \elapsed_time_ns_1_RNI0AND11_0_28\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__23465\,
            I => \N__23461\
        );

    \I__3464\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23458\
        );

    \I__3463\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23455\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__23458\,
            I => \N__23452\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__23455\,
            I => \N__23449\
        );

    \I__3460\ : Span4Mux_h
    port map (
            O => \N__23452\,
            I => \N__23446\
        );

    \I__3459\ : Span4Mux_h
    port map (
            O => \N__23449\,
            I => \N__23443\
        );

    \I__3458\ : Odrv4
    port map (
            O => \N__23446\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__23443\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__3456\ : InMux
    port map (
            O => \N__23438\,
            I => \N__23434\
        );

    \I__3455\ : InMux
    port map (
            O => \N__23437\,
            I => \N__23431\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__23434\,
            I => \N__23428\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__23431\,
            I => \elapsed_time_ns_1_RNIP3OD11_0_30\
        );

    \I__3452\ : Odrv4
    port map (
            O => \N__23428\,
            I => \elapsed_time_ns_1_RNIP3OD11_0_30\
        );

    \I__3451\ : InMux
    port map (
            O => \N__23423\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__3450\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23417\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__23417\,
            I => \N__23413\
        );

    \I__3448\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23408\
        );

    \I__3447\ : Span4Mux_v
    port map (
            O => \N__23413\,
            I => \N__23405\
        );

    \I__3446\ : InMux
    port map (
            O => \N__23412\,
            I => \N__23402\
        );

    \I__3445\ : InMux
    port map (
            O => \N__23411\,
            I => \N__23398\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__23408\,
            I => \N__23391\
        );

    \I__3443\ : Span4Mux_h
    port map (
            O => \N__23405\,
            I => \N__23391\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__23402\,
            I => \N__23391\
        );

    \I__3441\ : InMux
    port map (
            O => \N__23401\,
            I => \N__23388\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__23398\,
            I => \elapsed_time_ns_1_RNI40CED1_0_17\
        );

    \I__3439\ : Odrv4
    port map (
            O => \N__23391\,
            I => \elapsed_time_ns_1_RNI40CED1_0_17\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__23388\,
            I => \elapsed_time_ns_1_RNI40CED1_0_17\
        );

    \I__3437\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__23378\,
            I => \N__23372\
        );

    \I__3435\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23369\
        );

    \I__3434\ : InMux
    port map (
            O => \N__23376\,
            I => \N__23366\
        );

    \I__3433\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23363\
        );

    \I__3432\ : Span4Mux_h
    port map (
            O => \N__23372\,
            I => \N__23360\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__23369\,
            I => \N__23357\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__23366\,
            I => \N__23354\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__23363\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__23360\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__23357\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18\
        );

    \I__3426\ : Odrv4
    port map (
            O => \N__23354\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18\
        );

    \I__3425\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23342\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23337\
        );

    \I__3423\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23333\
        );

    \I__3422\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23330\
        );

    \I__3421\ : Span4Mux_v
    port map (
            O => \N__23337\,
            I => \N__23327\
        );

    \I__3420\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23324\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__23333\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__23330\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__23327\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__23324\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__23315\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3Z0Z_2_cascade_\
        );

    \I__3414\ : InMux
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__23309\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__3412\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__3410\ : Span4Mux_h
    port map (
            O => \N__23300\,
            I => \N__23296\
        );

    \I__3409\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23293\
        );

    \I__3408\ : Span4Mux_h
    port map (
            O => \N__23296\,
            I => \N__23288\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__23293\,
            I => \N__23288\
        );

    \I__3406\ : Odrv4
    port map (
            O => \N__23288\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__23285\,
            I => \N__23282\
        );

    \I__3404\ : InMux
    port map (
            O => \N__23282\,
            I => \N__23279\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23276\
        );

    \I__3402\ : Span4Mux_h
    port map (
            O => \N__23276\,
            I => \N__23272\
        );

    \I__3401\ : InMux
    port map (
            O => \N__23275\,
            I => \N__23269\
        );

    \I__3400\ : Span4Mux_v
    port map (
            O => \N__23272\,
            I => \N__23266\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__23269\,
            I => \N__23263\
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__23266\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__3397\ : Odrv12
    port map (
            O => \N__23263\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__3396\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23255\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__23255\,
            I => \elapsed_time_ns_1_RNI1BND11_0_29\
        );

    \I__3394\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23246\
        );

    \I__3393\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23246\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__23246\,
            I => \elapsed_time_ns_1_RNIP2ND11_0_21\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__23243\,
            I => \elapsed_time_ns_1_RNI1BND11_0_29_cascade_\
        );

    \I__3390\ : InMux
    port map (
            O => \N__23240\,
            I => \N__23237\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__23237\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_o5_0Z0Z_15\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__23234\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_o5_7Z0Z_15_cascade_\
        );

    \I__3387\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23228\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__23228\,
            I => \N__23225\
        );

    \I__3385\ : Span4Mux_h
    port map (
            O => \N__23225\,
            I => \N__23221\
        );

    \I__3384\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23218\
        );

    \I__3383\ : Span4Mux_h
    port map (
            O => \N__23221\,
            I => \N__23213\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__23218\,
            I => \N__23213\
        );

    \I__3381\ : Odrv4
    port map (
            O => \N__23213\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__3380\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23204\
        );

    \I__3379\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23204\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__23204\,
            I => \elapsed_time_ns_1_RNIO1ND11_0_20\
        );

    \I__3377\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23198\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__23198\,
            I => \N__23194\
        );

    \I__3375\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23191\
        );

    \I__3374\ : Span4Mux_h
    port map (
            O => \N__23194\,
            I => \N__23186\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__23191\,
            I => \N__23186\
        );

    \I__3372\ : Span4Mux_v
    port map (
            O => \N__23186\,
            I => \N__23183\
        );

    \I__3371\ : Odrv4
    port map (
            O => \N__23183\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__3370\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23174\
        );

    \I__3369\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23174\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__23174\,
            I => \elapsed_time_ns_1_RNIQ3ND11_0_22\
        );

    \I__3367\ : InMux
    port map (
            O => \N__23171\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__3366\ : InMux
    port map (
            O => \N__23168\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__3365\ : InMux
    port map (
            O => \N__23165\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__3364\ : InMux
    port map (
            O => \N__23162\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__3363\ : InMux
    port map (
            O => \N__23159\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__3362\ : InMux
    port map (
            O => \N__23156\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__3361\ : InMux
    port map (
            O => \N__23153\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__3360\ : InMux
    port map (
            O => \N__23150\,
            I => \bfn_9_15_0_\
        );

    \I__3359\ : InMux
    port map (
            O => \N__23147\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__3358\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23141\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__23141\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__3356\ : InMux
    port map (
            O => \N__23138\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__3355\ : InMux
    port map (
            O => \N__23135\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__3354\ : InMux
    port map (
            O => \N__23132\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__3353\ : InMux
    port map (
            O => \N__23129\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__3352\ : InMux
    port map (
            O => \N__23126\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__3351\ : InMux
    port map (
            O => \N__23123\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__3350\ : InMux
    port map (
            O => \N__23120\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__3349\ : InMux
    port map (
            O => \N__23117\,
            I => \bfn_9_14_0_\
        );

    \I__3348\ : IoInMux
    port map (
            O => \N__23114\,
            I => \N__23111\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__23111\,
            I => s4_phy_c
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__23108\,
            I => \N__23105\
        );

    \I__3345\ : InMux
    port map (
            O => \N__23105\,
            I => \N__23102\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__23102\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__23099\,
            I => \N__23096\
        );

    \I__3342\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23093\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__23093\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23087\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__23087\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__23084\,
            I => \N__23081\
        );

    \I__3337\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23078\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__23078\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__3335\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23072\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__23072\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__3333\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23066\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__23066\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__3331\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__23060\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__23057\,
            I => \N__23050\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__23056\,
            I => \N__23046\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__23055\,
            I => \N__23042\
        );

    \I__3326\ : InMux
    port map (
            O => \N__23054\,
            I => \N__23018\
        );

    \I__3325\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23018\
        );

    \I__3324\ : InMux
    port map (
            O => \N__23050\,
            I => \N__23018\
        );

    \I__3323\ : InMux
    port map (
            O => \N__23049\,
            I => \N__23018\
        );

    \I__3322\ : InMux
    port map (
            O => \N__23046\,
            I => \N__23018\
        );

    \I__3321\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23018\
        );

    \I__3320\ : InMux
    port map (
            O => \N__23042\,
            I => \N__23018\
        );

    \I__3319\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23018\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__23040\,
            I => \N__23014\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__23039\,
            I => \N__23010\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__23038\,
            I => \N__23006\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__23037\,
            I => \N__23002\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__23036\,
            I => \N__22999\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__23035\,
            I => \N__22995\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__23018\,
            I => \N__22991\
        );

    \I__3311\ : InMux
    port map (
            O => \N__23017\,
            I => \N__22974\
        );

    \I__3310\ : InMux
    port map (
            O => \N__23014\,
            I => \N__22974\
        );

    \I__3309\ : InMux
    port map (
            O => \N__23013\,
            I => \N__22974\
        );

    \I__3308\ : InMux
    port map (
            O => \N__23010\,
            I => \N__22974\
        );

    \I__3307\ : InMux
    port map (
            O => \N__23009\,
            I => \N__22974\
        );

    \I__3306\ : InMux
    port map (
            O => \N__23006\,
            I => \N__22974\
        );

    \I__3305\ : InMux
    port map (
            O => \N__23005\,
            I => \N__22974\
        );

    \I__3304\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22974\
        );

    \I__3303\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22965\
        );

    \I__3302\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22965\
        );

    \I__3301\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22965\
        );

    \I__3300\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22965\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__22991\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__22974\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__22965\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__22958\,
            I => \N__22955\
        );

    \I__3295\ : InMux
    port map (
            O => \N__22955\,
            I => \N__22950\
        );

    \I__3294\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22947\
        );

    \I__3293\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22944\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__22950\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__22947\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__22944\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__3289\ : InMux
    port map (
            O => \N__22937\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__3288\ : InMux
    port map (
            O => \N__22934\,
            I => \N__22929\
        );

    \I__3287\ : InMux
    port map (
            O => \N__22933\,
            I => \N__22924\
        );

    \I__3286\ : InMux
    port map (
            O => \N__22932\,
            I => \N__22924\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__22929\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__22924\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__3283\ : InMux
    port map (
            O => \N__22919\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__3282\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22911\
        );

    \I__3281\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22906\
        );

    \I__3280\ : InMux
    port map (
            O => \N__22914\,
            I => \N__22906\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__22911\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__22906\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__3277\ : InMux
    port map (
            O => \N__22901\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__22898\,
            I => \N__22894\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__22897\,
            I => \N__22891\
        );

    \I__3274\ : InMux
    port map (
            O => \N__22894\,
            I => \N__22887\
        );

    \I__3273\ : InMux
    port map (
            O => \N__22891\,
            I => \N__22884\
        );

    \I__3272\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22881\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__22887\,
            I => \N__22878\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__22884\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__22881\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__22878\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__3267\ : InMux
    port map (
            O => \N__22871\,
            I => \bfn_8_22_0_\
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__22868\,
            I => \N__22864\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__22867\,
            I => \N__22861\
        );

    \I__3264\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22857\
        );

    \I__3263\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22854\
        );

    \I__3262\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22851\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__22857\,
            I => \N__22848\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__22854\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__22851\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__22848\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__3257\ : InMux
    port map (
            O => \N__22841\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__22838\,
            I => \N__22835\
        );

    \I__3255\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22830\
        );

    \I__3254\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22827\
        );

    \I__3253\ : InMux
    port map (
            O => \N__22833\,
            I => \N__22824\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__22830\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__22827\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__22824\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__3249\ : InMux
    port map (
            O => \N__22817\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__22814\,
            I => \N__22811\
        );

    \I__3247\ : InMux
    port map (
            O => \N__22811\,
            I => \N__22806\
        );

    \I__3246\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22803\
        );

    \I__3245\ : InMux
    port map (
            O => \N__22809\,
            I => \N__22800\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__22806\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__22803\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__22800\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__3241\ : InMux
    port map (
            O => \N__22793\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__3240\ : InMux
    port map (
            O => \N__22790\,
            I => \N__22786\
        );

    \I__3239\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22783\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__22786\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__22783\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__3236\ : InMux
    port map (
            O => \N__22778\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__3235\ : InMux
    port map (
            O => \N__22775\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__3234\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22768\
        );

    \I__3233\ : InMux
    port map (
            O => \N__22771\,
            I => \N__22765\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__22768\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__22765\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__22760\,
            I => \N__22757\
        );

    \I__3229\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22752\
        );

    \I__3228\ : InMux
    port map (
            O => \N__22756\,
            I => \N__22749\
        );

    \I__3227\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22746\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__22752\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__22749\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__22746\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__3223\ : InMux
    port map (
            O => \N__22739\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__3222\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22731\
        );

    \I__3221\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22726\
        );

    \I__3220\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22726\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__22731\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__22726\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__3217\ : InMux
    port map (
            O => \N__22721\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__3216\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22713\
        );

    \I__3215\ : InMux
    port map (
            O => \N__22717\,
            I => \N__22708\
        );

    \I__3214\ : InMux
    port map (
            O => \N__22716\,
            I => \N__22708\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__22713\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__22708\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__3211\ : InMux
    port map (
            O => \N__22703\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__3210\ : CascadeMux
    port map (
            O => \N__22700\,
            I => \N__22696\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__22699\,
            I => \N__22693\
        );

    \I__3208\ : InMux
    port map (
            O => \N__22696\,
            I => \N__22689\
        );

    \I__3207\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22686\
        );

    \I__3206\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22683\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__22689\,
            I => \N__22680\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__22686\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__22683\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__22680\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__3201\ : InMux
    port map (
            O => \N__22673\,
            I => \bfn_8_21_0_\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__22670\,
            I => \N__22666\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__22669\,
            I => \N__22663\
        );

    \I__3198\ : InMux
    port map (
            O => \N__22666\,
            I => \N__22659\
        );

    \I__3197\ : InMux
    port map (
            O => \N__22663\,
            I => \N__22656\
        );

    \I__3196\ : InMux
    port map (
            O => \N__22662\,
            I => \N__22653\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__22659\,
            I => \N__22650\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__22656\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__22653\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__22650\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__3191\ : InMux
    port map (
            O => \N__22643\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__22640\,
            I => \N__22637\
        );

    \I__3189\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22632\
        );

    \I__3188\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22629\
        );

    \I__3187\ : InMux
    port map (
            O => \N__22635\,
            I => \N__22626\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__22632\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__22629\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__22626\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__3183\ : InMux
    port map (
            O => \N__22619\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__22616\,
            I => \N__22613\
        );

    \I__3181\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22608\
        );

    \I__3180\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22605\
        );

    \I__3179\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22602\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__22608\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__22605\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__22602\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__3175\ : InMux
    port map (
            O => \N__22595\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__22592\,
            I => \N__22589\
        );

    \I__3173\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22584\
        );

    \I__3172\ : InMux
    port map (
            O => \N__22588\,
            I => \N__22581\
        );

    \I__3171\ : InMux
    port map (
            O => \N__22587\,
            I => \N__22578\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__22584\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__22581\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__22578\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__3167\ : InMux
    port map (
            O => \N__22571\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__3165\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22560\
        );

    \I__3164\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22557\
        );

    \I__3163\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22554\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__22560\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__22557\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__22554\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__3159\ : InMux
    port map (
            O => \N__22547\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__3158\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22539\
        );

    \I__3157\ : InMux
    port map (
            O => \N__22543\,
            I => \N__22534\
        );

    \I__3156\ : InMux
    port map (
            O => \N__22542\,
            I => \N__22534\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__22539\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__22534\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__3153\ : InMux
    port map (
            O => \N__22529\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__3152\ : InMux
    port map (
            O => \N__22526\,
            I => \N__22521\
        );

    \I__3151\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22516\
        );

    \I__3150\ : InMux
    port map (
            O => \N__22524\,
            I => \N__22516\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__22521\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__22516\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__3147\ : InMux
    port map (
            O => \N__22511\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__22508\,
            I => \N__22505\
        );

    \I__3145\ : InMux
    port map (
            O => \N__22505\,
            I => \N__22501\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__22504\,
            I => \N__22498\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__22501\,
            I => \N__22494\
        );

    \I__3142\ : InMux
    port map (
            O => \N__22498\,
            I => \N__22491\
        );

    \I__3141\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22488\
        );

    \I__3140\ : Span4Mux_h
    port map (
            O => \N__22494\,
            I => \N__22485\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__22491\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__22488\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__22485\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__3136\ : InMux
    port map (
            O => \N__22478\,
            I => \bfn_8_20_0_\
        );

    \I__3135\ : CascadeMux
    port map (
            O => \N__22475\,
            I => \N__22471\
        );

    \I__3134\ : CascadeMux
    port map (
            O => \N__22474\,
            I => \N__22468\
        );

    \I__3133\ : InMux
    port map (
            O => \N__22471\,
            I => \N__22464\
        );

    \I__3132\ : InMux
    port map (
            O => \N__22468\,
            I => \N__22461\
        );

    \I__3131\ : InMux
    port map (
            O => \N__22467\,
            I => \N__22458\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__22464\,
            I => \N__22455\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__22461\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__22458\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__22455\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__3126\ : InMux
    port map (
            O => \N__22448\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__22445\,
            I => \N__22442\
        );

    \I__3124\ : InMux
    port map (
            O => \N__22442\,
            I => \N__22437\
        );

    \I__3123\ : InMux
    port map (
            O => \N__22441\,
            I => \N__22434\
        );

    \I__3122\ : InMux
    port map (
            O => \N__22440\,
            I => \N__22431\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__22437\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__22434\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__22431\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__3118\ : InMux
    port map (
            O => \N__22424\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__22421\,
            I => \N__22418\
        );

    \I__3116\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22413\
        );

    \I__3115\ : InMux
    port map (
            O => \N__22417\,
            I => \N__22410\
        );

    \I__3114\ : InMux
    port map (
            O => \N__22416\,
            I => \N__22407\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__22413\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__22410\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__22407\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__3110\ : InMux
    port map (
            O => \N__22400\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__3108\ : InMux
    port map (
            O => \N__22394\,
            I => \N__22389\
        );

    \I__3107\ : InMux
    port map (
            O => \N__22393\,
            I => \N__22386\
        );

    \I__3106\ : InMux
    port map (
            O => \N__22392\,
            I => \N__22383\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__22389\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__22386\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__22383\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__3102\ : InMux
    port map (
            O => \N__22376\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__3101\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22369\
        );

    \I__3100\ : InMux
    port map (
            O => \N__22372\,
            I => \N__22366\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__22369\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__22366\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__3097\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22358\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__22358\,
            I => \N__22354\
        );

    \I__3095\ : InMux
    port map (
            O => \N__22357\,
            I => \N__22351\
        );

    \I__3094\ : Odrv4
    port map (
            O => \N__22354\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__22351\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__3092\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__22343\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16\
        );

    \I__3090\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22335\
        );

    \I__3089\ : InMux
    port map (
            O => \N__22339\,
            I => \N__22330\
        );

    \I__3088\ : InMux
    port map (
            O => \N__22338\,
            I => \N__22330\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__22335\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__22330\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__22325\,
            I => \N__22321\
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__22324\,
            I => \N__22318\
        );

    \I__3083\ : InMux
    port map (
            O => \N__22321\,
            I => \N__22314\
        );

    \I__3082\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22309\
        );

    \I__3081\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22309\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__22314\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__22309\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\
        );

    \I__3078\ : InMux
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__22301\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15\
        );

    \I__3076\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__22295\,
            I => \N__22291\
        );

    \I__3074\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22288\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__22291\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__22288\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__22283\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__3069\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22273\
        );

    \I__3068\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22270\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__22273\,
            I => \N__22266\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22263\
        );

    \I__3065\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22260\
        );

    \I__3064\ : Odrv4
    port map (
            O => \N__22266\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__22263\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__22260\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\
        );

    \I__3061\ : InMux
    port map (
            O => \N__22253\,
            I => \bfn_8_19_0_\
        );

    \I__3060\ : InMux
    port map (
            O => \N__22250\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__22247\,
            I => \N__22244\
        );

    \I__3058\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22239\
        );

    \I__3057\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22236\
        );

    \I__3056\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22233\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__22239\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__22236\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__22233\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__3052\ : InMux
    port map (
            O => \N__22226\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__3050\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22215\
        );

    \I__3049\ : InMux
    port map (
            O => \N__22219\,
            I => \N__22212\
        );

    \I__3048\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22209\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__22215\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__22212\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__22209\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__3044\ : InMux
    port map (
            O => \N__22202\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__22199\,
            I => \N__22196\
        );

    \I__3042\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22191\
        );

    \I__3041\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22188\
        );

    \I__3040\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22185\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__22191\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__22188\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__22185\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__3036\ : InMux
    port map (
            O => \N__22178\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__3035\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__22172\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31\
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__3032\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__22163\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5\
        );

    \I__3030\ : InMux
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__22157\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__22154\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_\
        );

    \I__3027\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22147\
        );

    \I__3026\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22144\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__22147\,
            I => \N__22141\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__22144\,
            I => \N__22138\
        );

    \I__3023\ : Span4Mux_v
    port map (
            O => \N__22141\,
            I => \N__22134\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__22138\,
            I => \N__22131\
        );

    \I__3021\ : InMux
    port map (
            O => \N__22137\,
            I => \N__22128\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__22134\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__22131\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__22128\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__3017\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22115\
        );

    \I__3016\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22115\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__22115\,
            I => \N__22111\
        );

    \I__3014\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22108\
        );

    \I__3013\ : Span4Mux_v
    port map (
            O => \N__22111\,
            I => \N__22105\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__22108\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__22105\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__3010\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22095\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__22099\,
            I => \N__22092\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__22098\,
            I => \N__22089\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__22095\,
            I => \N__22086\
        );

    \I__3006\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22083\
        );

    \I__3005\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22080\
        );

    \I__3004\ : Span4Mux_v
    port map (
            O => \N__22086\,
            I => \N__22075\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__22083\,
            I => \N__22075\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__22080\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__22075\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__3000\ : InMux
    port map (
            O => \N__22070\,
            I => \N__22066\
        );

    \I__2999\ : InMux
    port map (
            O => \N__22069\,
            I => \N__22062\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__22066\,
            I => \N__22058\
        );

    \I__2997\ : InMux
    port map (
            O => \N__22065\,
            I => \N__22055\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__22062\,
            I => \N__22052\
        );

    \I__2995\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22049\
        );

    \I__2994\ : Odrv12
    port map (
            O => \N__22058\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__22055\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__22052\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__22049\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__2990\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22037\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__22037\,
            I => \N__22031\
        );

    \I__2988\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22028\
        );

    \I__2987\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22025\
        );

    \I__2986\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22022\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__22031\,
            I => \N__22015\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__22028\,
            I => \N__22015\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__22025\,
            I => \N__22015\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__22022\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__22015\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__22010\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__22007\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__22004\,
            I => \N__22000\
        );

    \I__2977\ : InMux
    port map (
            O => \N__22003\,
            I => \N__21997\
        );

    \I__2976\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21994\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__21997\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__21994\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__21989\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_\
        );

    \I__2972\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21983\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__21983\,
            I => \N__21980\
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__21980\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__21977\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_\
        );

    \I__2968\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__21971\,
            I => \N__21968\
        );

    \I__2966\ : Odrv12
    port map (
            O => \N__21968\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17\
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__21965\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__21962\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31_cascade_\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__21959\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31_cascade_\
        );

    \I__2962\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21953\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__21953\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2\
        );

    \I__2960\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__2958\ : Span4Mux_v
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__21941\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__2955\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21931\
        );

    \I__2954\ : InMux
    port map (
            O => \N__21934\,
            I => \N__21926\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__21931\,
            I => \N__21923\
        );

    \I__2952\ : InMux
    port map (
            O => \N__21930\,
            I => \N__21917\
        );

    \I__2951\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21917\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__21926\,
            I => \N__21912\
        );

    \I__2949\ : Span12Mux_s8_h
    port map (
            O => \N__21923\,
            I => \N__21912\
        );

    \I__2948\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21909\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__21917\,
            I => \N__21906\
        );

    \I__2946\ : Odrv12
    port map (
            O => \N__21912\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__21909\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__21906\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__21899\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14_cascade_\
        );

    \I__2942\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21892\
        );

    \I__2941\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21889\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__21892\,
            I => \N__21882\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__21889\,
            I => \N__21882\
        );

    \I__2938\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21879\
        );

    \I__2937\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21876\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__21882\,
            I => \elapsed_time_ns_1_RNIL13KD1_0_9\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__21879\,
            I => \elapsed_time_ns_1_RNIL13KD1_0_9\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__21876\,
            I => \elapsed_time_ns_1_RNIL13KD1_0_9\
        );

    \I__2933\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21865\
        );

    \I__2932\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21862\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__21865\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_1Z0Z_9\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__21862\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_1Z0Z_9\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__21857\,
            I => \N__21853\
        );

    \I__2928\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21850\
        );

    \I__2927\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21846\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__21850\,
            I => \N__21843\
        );

    \I__2925\ : InMux
    port map (
            O => \N__21849\,
            I => \N__21840\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__21846\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__21843\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__21840\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__21833\,
            I => \N__21827\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__21832\,
            I => \N__21820\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__21831\,
            I => \N__21817\
        );

    \I__2918\ : InMux
    port map (
            O => \N__21830\,
            I => \N__21811\
        );

    \I__2917\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21811\
        );

    \I__2916\ : InMux
    port map (
            O => \N__21826\,
            I => \N__21806\
        );

    \I__2915\ : InMux
    port map (
            O => \N__21825\,
            I => \N__21806\
        );

    \I__2914\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21801\
        );

    \I__2913\ : InMux
    port map (
            O => \N__21823\,
            I => \N__21801\
        );

    \I__2912\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21796\
        );

    \I__2911\ : InMux
    port map (
            O => \N__21817\,
            I => \N__21796\
        );

    \I__2910\ : InMux
    port map (
            O => \N__21816\,
            I => \N__21793\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__21811\,
            I => \phase_controller_inst1.stoper_hc.N_315\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__21806\,
            I => \phase_controller_inst1.stoper_hc.N_315\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__21801\,
            I => \phase_controller_inst1.stoper_hc.N_315\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__21796\,
            I => \phase_controller_inst1.stoper_hc.N_315\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__21793\,
            I => \phase_controller_inst1.stoper_hc.N_315\
        );

    \I__2904\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21778\
        );

    \I__2903\ : InMux
    port map (
            O => \N__21781\,
            I => \N__21773\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__21778\,
            I => \N__21770\
        );

    \I__2901\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21765\
        );

    \I__2900\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21765\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__21773\,
            I => \elapsed_time_ns_1_RNIO0MD11_0_11\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__21770\,
            I => \elapsed_time_ns_1_RNIO0MD11_0_11\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__21765\,
            I => \elapsed_time_ns_1_RNIO0MD11_0_11\
        );

    \I__2896\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21754\
        );

    \I__2895\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21751\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__21754\,
            I => \elapsed_time_ns_1_RNIR4ND11_0_23\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__21751\,
            I => \elapsed_time_ns_1_RNIR4ND11_0_23\
        );

    \I__2892\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21742\
        );

    \I__2891\ : InMux
    port map (
            O => \N__21745\,
            I => \N__21739\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__21742\,
            I => \N__21734\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__21739\,
            I => \N__21734\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__21734\,
            I => \elapsed_time_ns_1_RNIS5ND11_0_24\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__2886\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21724\
        );

    \I__2885\ : CascadeMux
    port map (
            O => \N__21727\,
            I => \N__21721\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__21724\,
            I => \N__21718\
        );

    \I__2883\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21715\
        );

    \I__2882\ : Span4Mux_h
    port map (
            O => \N__21718\,
            I => \N__21712\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__21715\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__21712\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2879\ : InMux
    port map (
            O => \N__21707\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2878\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__21701\,
            I => \N__21697\
        );

    \I__2876\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21694\
        );

    \I__2875\ : Span4Mux_v
    port map (
            O => \N__21697\,
            I => \N__21691\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__21694\,
            I => \N__21688\
        );

    \I__2873\ : Odrv4
    port map (
            O => \N__21691\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__21688\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2871\ : InMux
    port map (
            O => \N__21683\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2870\ : InMux
    port map (
            O => \N__21680\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2869\ : InMux
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__21674\,
            I => \N__21667\
        );

    \I__2867\ : InMux
    port map (
            O => \N__21673\,
            I => \N__21664\
        );

    \I__2866\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21656\
        );

    \I__2865\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21656\
        );

    \I__2864\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21653\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__21667\,
            I => \N__21646\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__21664\,
            I => \N__21646\
        );

    \I__2861\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21643\
        );

    \I__2860\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21638\
        );

    \I__2859\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21638\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__21656\,
            I => \N__21635\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__21653\,
            I => \N__21632\
        );

    \I__2856\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21627\
        );

    \I__2855\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21627\
        );

    \I__2854\ : Span4Mux_v
    port map (
            O => \N__21646\,
            I => \N__21624\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__21643\,
            I => \N__21619\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__21638\,
            I => \N__21619\
        );

    \I__2851\ : Span4Mux_v
    port map (
            O => \N__21635\,
            I => \N__21616\
        );

    \I__2850\ : Span12Mux_s8_h
    port map (
            O => \N__21632\,
            I => \N__21613\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__21627\,
            I => \N__21610\
        );

    \I__2848\ : Span4Mux_h
    port map (
            O => \N__21624\,
            I => \N__21605\
        );

    \I__2847\ : Span4Mux_v
    port map (
            O => \N__21619\,
            I => \N__21605\
        );

    \I__2846\ : Span4Mux_h
    port map (
            O => \N__21616\,
            I => \N__21602\
        );

    \I__2845\ : Odrv12
    port map (
            O => \N__21613\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2844\ : Odrv12
    port map (
            O => \N__21610\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__21605\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__21602\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2841\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21590\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__21590\,
            I => \N__21586\
        );

    \I__2839\ : InMux
    port map (
            O => \N__21589\,
            I => \N__21583\
        );

    \I__2838\ : Odrv12
    port map (
            O => \N__21586\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_14\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__21583\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_14\
        );

    \I__2836\ : InMux
    port map (
            O => \N__21578\,
            I => \N__21572\
        );

    \I__2835\ : InMux
    port map (
            O => \N__21577\,
            I => \N__21572\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__21572\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2833\ : InMux
    port map (
            O => \N__21569\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__21566\,
            I => \N__21563\
        );

    \I__2831\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21560\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__21560\,
            I => \N__21556\
        );

    \I__2829\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21553\
        );

    \I__2828\ : Odrv12
    port map (
            O => \N__21556\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__21553\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2826\ : InMux
    port map (
            O => \N__21548\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2825\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21542\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__21542\,
            I => \N__21538\
        );

    \I__2823\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21535\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__21538\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__21535\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2820\ : InMux
    port map (
            O => \N__21530\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2819\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21521\
        );

    \I__2818\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21521\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__21521\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2816\ : InMux
    port map (
            O => \N__21518\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__21515\,
            I => \N__21512\
        );

    \I__2814\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21508\
        );

    \I__2813\ : InMux
    port map (
            O => \N__21511\,
            I => \N__21505\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__21508\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__21505\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2810\ : InMux
    port map (
            O => \N__21500\,
            I => \bfn_8_13_0_\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__21497\,
            I => \N__21494\
        );

    \I__2808\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21488\
        );

    \I__2807\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21488\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__21488\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2805\ : InMux
    port map (
            O => \N__21485\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2804\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21475\
        );

    \I__2802\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21472\
        );

    \I__2801\ : Span4Mux_h
    port map (
            O => \N__21475\,
            I => \N__21469\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__21472\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__21469\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2798\ : InMux
    port map (
            O => \N__21464\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2797\ : InMux
    port map (
            O => \N__21461\,
            I => \N__21457\
        );

    \I__2796\ : InMux
    port map (
            O => \N__21460\,
            I => \N__21454\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__21457\,
            I => \N__21451\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__21454\,
            I => \N__21448\
        );

    \I__2793\ : Span4Mux_h
    port map (
            O => \N__21451\,
            I => \N__21445\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__21448\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2791\ : Odrv4
    port map (
            O => \N__21445\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2790\ : InMux
    port map (
            O => \N__21440\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2789\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21434\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__21434\,
            I => \N__21431\
        );

    \I__2787\ : Span4Mux_v
    port map (
            O => \N__21431\,
            I => \N__21427\
        );

    \I__2786\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21424\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__21427\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__21424\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2783\ : InMux
    port map (
            O => \N__21419\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__21416\,
            I => \N__21413\
        );

    \I__2781\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21410\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__21410\,
            I => \N__21406\
        );

    \I__2779\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21403\
        );

    \I__2778\ : Odrv12
    port map (
            O => \N__21406\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__21403\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2776\ : InMux
    port map (
            O => \N__21398\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2775\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21389\
        );

    \I__2774\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21389\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__21389\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2772\ : InMux
    port map (
            O => \N__21386\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__21383\,
            I => \N__21379\
        );

    \I__2770\ : InMux
    port map (
            O => \N__21382\,
            I => \N__21376\
        );

    \I__2769\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21373\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__21376\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__21373\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2766\ : InMux
    port map (
            O => \N__21368\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2765\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21362\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__21362\,
            I => \N__21359\
        );

    \I__2763\ : Span4Mux_h
    port map (
            O => \N__21359\,
            I => \N__21355\
        );

    \I__2762\ : InMux
    port map (
            O => \N__21358\,
            I => \N__21352\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__21355\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__21352\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2759\ : InMux
    port map (
            O => \N__21347\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__21344\,
            I => \N__21341\
        );

    \I__2757\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21338\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__21338\,
            I => \N__21334\
        );

    \I__2755\ : InMux
    port map (
            O => \N__21337\,
            I => \N__21331\
        );

    \I__2754\ : Odrv12
    port map (
            O => \N__21334\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__21331\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2752\ : InMux
    port map (
            O => \N__21326\,
            I => \bfn_8_12_0_\
        );

    \I__2751\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21317\
        );

    \I__2750\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21317\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__21317\,
            I => \N__21314\
        );

    \I__2748\ : Odrv12
    port map (
            O => \N__21314\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2747\ : InMux
    port map (
            O => \N__21311\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__21308\,
            I => \N__21305\
        );

    \I__2745\ : InMux
    port map (
            O => \N__21305\,
            I => \N__21299\
        );

    \I__2744\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21299\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__21299\,
            I => \N__21296\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__21296\,
            I => \N__21293\
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__21293\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2740\ : InMux
    port map (
            O => \N__21290\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2739\ : InMux
    port map (
            O => \N__21287\,
            I => \N__21281\
        );

    \I__2738\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21281\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__21281\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2736\ : InMux
    port map (
            O => \N__21278\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__21275\,
            I => \N__21271\
        );

    \I__2734\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21268\
        );

    \I__2733\ : InMux
    port map (
            O => \N__21271\,
            I => \N__21265\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__21268\,
            I => \N__21262\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__21265\,
            I => \N__21259\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__21262\,
            I => \N__21256\
        );

    \I__2729\ : Span12Mux_v
    port map (
            O => \N__21259\,
            I => \N__21250\
        );

    \I__2728\ : Sp12to4
    port map (
            O => \N__21256\,
            I => \N__21250\
        );

    \I__2727\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21247\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__21250\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__21247\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2724\ : InMux
    port map (
            O => \N__21242\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2723\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21235\
        );

    \I__2722\ : InMux
    port map (
            O => \N__21238\,
            I => \N__21231\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__21235\,
            I => \N__21228\
        );

    \I__2720\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21225\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__21231\,
            I => \N__21220\
        );

    \I__2718\ : Span4Mux_h
    port map (
            O => \N__21228\,
            I => \N__21220\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__21225\,
            I => \N__21216\
        );

    \I__2716\ : Span4Mux_h
    port map (
            O => \N__21220\,
            I => \N__21213\
        );

    \I__2715\ : InMux
    port map (
            O => \N__21219\,
            I => \N__21210\
        );

    \I__2714\ : Odrv12
    port map (
            O => \N__21216\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__21213\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__21210\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2711\ : InMux
    port map (
            O => \N__21203\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__21200\,
            I => \N__21197\
        );

    \I__2709\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21194\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__21194\,
            I => \N__21189\
        );

    \I__2707\ : InMux
    port map (
            O => \N__21193\,
            I => \N__21186\
        );

    \I__2706\ : InMux
    port map (
            O => \N__21192\,
            I => \N__21183\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__21189\,
            I => \N__21180\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__21186\,
            I => \N__21175\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__21183\,
            I => \N__21175\
        );

    \I__2702\ : Span4Mux_h
    port map (
            O => \N__21180\,
            I => \N__21170\
        );

    \I__2701\ : Span4Mux_v
    port map (
            O => \N__21175\,
            I => \N__21170\
        );

    \I__2700\ : Odrv4
    port map (
            O => \N__21170\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2699\ : InMux
    port map (
            O => \N__21167\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__21164\,
            I => \N__21161\
        );

    \I__2697\ : InMux
    port map (
            O => \N__21161\,
            I => \N__21158\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__21158\,
            I => \N__21154\
        );

    \I__2695\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21151\
        );

    \I__2694\ : Span4Mux_h
    port map (
            O => \N__21154\,
            I => \N__21145\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__21151\,
            I => \N__21145\
        );

    \I__2692\ : InMux
    port map (
            O => \N__21150\,
            I => \N__21142\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__21145\,
            I => \N__21137\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__21142\,
            I => \N__21137\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__21137\,
            I => \N__21134\
        );

    \I__2688\ : Odrv4
    port map (
            O => \N__21134\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2687\ : InMux
    port map (
            O => \N__21131\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__21128\,
            I => \N__21123\
        );

    \I__2685\ : InMux
    port map (
            O => \N__21127\,
            I => \N__21120\
        );

    \I__2684\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21117\
        );

    \I__2683\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21114\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__21120\,
            I => \N__21109\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__21117\,
            I => \N__21109\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__21114\,
            I => \N__21106\
        );

    \I__2679\ : Span4Mux_v
    port map (
            O => \N__21109\,
            I => \N__21103\
        );

    \I__2678\ : Odrv12
    port map (
            O => \N__21106\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2677\ : Odrv4
    port map (
            O => \N__21103\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2676\ : InMux
    port map (
            O => \N__21098\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__21095\,
            I => \N__21092\
        );

    \I__2674\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21088\
        );

    \I__2673\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21085\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__21088\,
            I => \N__21081\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__21085\,
            I => \N__21078\
        );

    \I__2670\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21075\
        );

    \I__2669\ : Span4Mux_h
    port map (
            O => \N__21081\,
            I => \N__21072\
        );

    \I__2668\ : Span4Mux_v
    port map (
            O => \N__21078\,
            I => \N__21067\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__21075\,
            I => \N__21067\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__21072\,
            I => \N__21064\
        );

    \I__2665\ : Span4Mux_h
    port map (
            O => \N__21067\,
            I => \N__21061\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__21064\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__21061\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2662\ : InMux
    port map (
            O => \N__21056\,
            I => \bfn_8_11_0_\
        );

    \I__2661\ : InMux
    port map (
            O => \N__21053\,
            I => \N__21050\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__21050\,
            I => \N__21045\
        );

    \I__2659\ : InMux
    port map (
            O => \N__21049\,
            I => \N__21042\
        );

    \I__2658\ : InMux
    port map (
            O => \N__21048\,
            I => \N__21039\
        );

    \I__2657\ : Span4Mux_h
    port map (
            O => \N__21045\,
            I => \N__21034\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__21042\,
            I => \N__21034\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__21039\,
            I => \N__21031\
        );

    \I__2654\ : Span4Mux_h
    port map (
            O => \N__21034\,
            I => \N__21028\
        );

    \I__2653\ : Odrv12
    port map (
            O => \N__21031\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__21028\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2651\ : InMux
    port map (
            O => \N__21023\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2650\ : InMux
    port map (
            O => \N__21020\,
            I => \N__21014\
        );

    \I__2649\ : InMux
    port map (
            O => \N__21019\,
            I => \N__21014\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__21014\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2647\ : InMux
    port map (
            O => \N__21011\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2646\ : InMux
    port map (
            O => \N__21008\,
            I => \N__21005\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__21005\,
            I => \N__21001\
        );

    \I__2644\ : InMux
    port map (
            O => \N__21004\,
            I => \N__20998\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__21001\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__20998\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2641\ : InMux
    port map (
            O => \N__20993\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2640\ : InMux
    port map (
            O => \N__20990\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__2639\ : InMux
    port map (
            O => \N__20987\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__2638\ : InMux
    port map (
            O => \N__20984\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__2637\ : InMux
    port map (
            O => \N__20981\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__2636\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20975\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20972\
        );

    \I__2634\ : Span4Mux_h
    port map (
            O => \N__20972\,
            I => \N__20969\
        );

    \I__2633\ : Span4Mux_v
    port map (
            O => \N__20969\,
            I => \N__20966\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__20966\,
            I => il_min_comp2_c
        );

    \I__2631\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__20960\,
            I => \N__20957\
        );

    \I__2629\ : Span4Mux_h
    port map (
            O => \N__20957\,
            I => \N__20954\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__20951\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2626\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20945\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__20945\,
            I => \N__20942\
        );

    \I__2624\ : Span4Mux_h
    port map (
            O => \N__20942\,
            I => \N__20939\
        );

    \I__2623\ : Span4Mux_h
    port map (
            O => \N__20939\,
            I => \N__20936\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__20936\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2621\ : InMux
    port map (
            O => \N__20933\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__2619\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20924\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__20924\,
            I => \N__20921\
        );

    \I__2617\ : Span12Mux_s8_h
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__2616\ : Odrv12
    port map (
            O => \N__20918\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2615\ : InMux
    port map (
            O => \N__20915\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2614\ : InMux
    port map (
            O => \N__20912\,
            I => \bfn_7_20_0_\
        );

    \I__2613\ : InMux
    port map (
            O => \N__20909\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__2612\ : InMux
    port map (
            O => \N__20906\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__2611\ : InMux
    port map (
            O => \N__20903\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__2609\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__20894\,
            I => \N__20890\
        );

    \I__2607\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20887\
        );

    \I__2606\ : Span4Mux_v
    port map (
            O => \N__20890\,
            I => \N__20882\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__20887\,
            I => \N__20882\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__20882\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__2603\ : InMux
    port map (
            O => \N__20879\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__2602\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20873\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__20873\,
            I => \N__20869\
        );

    \I__2600\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20866\
        );

    \I__2599\ : Span4Mux_h
    port map (
            O => \N__20869\,
            I => \N__20861\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20861\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__20861\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__2596\ : InMux
    port map (
            O => \N__20858\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__2595\ : InMux
    port map (
            O => \N__20855\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__2594\ : InMux
    port map (
            O => \N__20852\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__2593\ : InMux
    port map (
            O => \N__20849\,
            I => \bfn_7_21_0_\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__20846\,
            I => \N__20843\
        );

    \I__2591\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20840\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__20840\,
            I => \N__20836\
        );

    \I__2589\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20833\
        );

    \I__2588\ : Odrv12
    port map (
            O => \N__20836\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__20833\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__2586\ : InMux
    port map (
            O => \N__20828\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__20825\,
            I => \N__20822\
        );

    \I__2584\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20819\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__20819\,
            I => \N__20815\
        );

    \I__2582\ : InMux
    port map (
            O => \N__20818\,
            I => \N__20812\
        );

    \I__2581\ : Span4Mux_h
    port map (
            O => \N__20815\,
            I => \N__20809\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__20812\,
            I => \N__20806\
        );

    \I__2579\ : Odrv4
    port map (
            O => \N__20809\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__20806\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__2577\ : InMux
    port map (
            O => \N__20801\,
            I => \bfn_7_19_0_\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__20798\,
            I => \N__20795\
        );

    \I__2575\ : InMux
    port map (
            O => \N__20795\,
            I => \N__20791\
        );

    \I__2574\ : InMux
    port map (
            O => \N__20794\,
            I => \N__20788\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__20791\,
            I => \N__20785\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__20788\,
            I => \N__20782\
        );

    \I__2571\ : Odrv12
    port map (
            O => \N__20785\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__20782\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__2569\ : InMux
    port map (
            O => \N__20777\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__20774\,
            I => \N__20770\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__20773\,
            I => \N__20767\
        );

    \I__2566\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20764\
        );

    \I__2565\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20761\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20758\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__20761\,
            I => \N__20755\
        );

    \I__2562\ : Odrv12
    port map (
            O => \N__20758\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__20755\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__2560\ : InMux
    port map (
            O => \N__20750\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__2559\ : InMux
    port map (
            O => \N__20747\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__20744\,
            I => \N__20741\
        );

    \I__2557\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20736\
        );

    \I__2556\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20731\
        );

    \I__2555\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20731\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__20736\,
            I => \N__20726\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__20731\,
            I => \N__20726\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__20726\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\
        );

    \I__2551\ : InMux
    port map (
            O => \N__20723\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__2550\ : InMux
    port map (
            O => \N__20720\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__2549\ : InMux
    port map (
            O => \N__20717\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__2548\ : InMux
    port map (
            O => \N__20714\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__2547\ : InMux
    port map (
            O => \N__20711\,
            I => \N__20708\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__20708\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__20705\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_\
        );

    \I__2544\ : InMux
    port map (
            O => \N__20702\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__2543\ : InMux
    port map (
            O => \N__20699\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__2542\ : InMux
    port map (
            O => \N__20696\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__2541\ : InMux
    port map (
            O => \N__20693\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__2540\ : InMux
    port map (
            O => \N__20690\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__2539\ : InMux
    port map (
            O => \N__20687\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__2538\ : InMux
    port map (
            O => \N__20684\,
            I => \N__20681\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__20681\,
            I => \N__20678\
        );

    \I__2536\ : Odrv12
    port map (
            O => \N__20678\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__20675\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__20672\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4_cascade_\
        );

    \I__2533\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20666\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__20666\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__20663\,
            I => \elapsed_time_ns_1_RNIP1MD11_0_12_cascade_\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__20660\,
            I => \N__20657\
        );

    \I__2529\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20654\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__20654\,
            I => \N__20649\
        );

    \I__2527\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20644\
        );

    \I__2526\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20644\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__20649\,
            I => \elapsed_time_ns_1_RNIP1MD11_0_12\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__20644\,
            I => \elapsed_time_ns_1_RNIP1MD11_0_12\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__20639\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10_cascade_\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__20636\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2_cascade_\
        );

    \I__2521\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20629\
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__20632\,
            I => \N__20625\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__20629\,
            I => \N__20621\
        );

    \I__2518\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20614\
        );

    \I__2517\ : InMux
    port map (
            O => \N__20625\,
            I => \N__20614\
        );

    \I__2516\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20614\
        );

    \I__2515\ : Odrv4
    port map (
            O => \N__20621\,
            I => \elapsed_time_ns_1_RNIQ2MD11_0_13\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__20614\,
            I => \elapsed_time_ns_1_RNIQ2MD11_0_13\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__20609\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18_cascade_\
        );

    \I__2512\ : InMux
    port map (
            O => \N__20606\,
            I => \N__20603\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__20603\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__20600\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__20597\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16_cascade_\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__20594\,
            I => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9_cascade_\
        );

    \I__2507\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20588\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__20588\,
            I => \N__20585\
        );

    \I__2505\ : Span4Mux_h
    port map (
            O => \N__20585\,
            I => \N__20582\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__20582\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__20579\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\
        );

    \I__2502\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20573\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__20573\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\
        );

    \I__2500\ : InMux
    port map (
            O => \N__20570\,
            I => \N__20567\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__20567\,
            I => \N__20564\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__20564\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2497\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20558\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__20558\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2495\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20549\
        );

    \I__2494\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20541\
        );

    \I__2493\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20541\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__20552\,
            I => \N__20538\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__20549\,
            I => \N__20535\
        );

    \I__2490\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20531\
        );

    \I__2489\ : InMux
    port map (
            O => \N__20547\,
            I => \N__20526\
        );

    \I__2488\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20526\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__20541\,
            I => \N__20522\
        );

    \I__2486\ : InMux
    port map (
            O => \N__20538\,
            I => \N__20519\
        );

    \I__2485\ : Span4Mux_s3_h
    port map (
            O => \N__20535\,
            I => \N__20516\
        );

    \I__2484\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20513\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__20531\,
            I => \N__20510\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__20526\,
            I => \N__20507\
        );

    \I__2481\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20504\
        );

    \I__2480\ : Span4Mux_v
    port map (
            O => \N__20522\,
            I => \N__20499\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__20519\,
            I => \N__20499\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__20516\,
            I => \N__20494\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__20513\,
            I => \N__20494\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__20510\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2475\ : Odrv12
    port map (
            O => \N__20507\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__20504\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__20499\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2472\ : Odrv4
    port map (
            O => \N__20494\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2471\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20480\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__20480\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\
        );

    \I__2469\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20474\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__20474\,
            I => \N__20471\
        );

    \I__2467\ : Span12Mux_v
    port map (
            O => \N__20471\,
            I => \N__20468\
        );

    \I__2466\ : Odrv12
    port map (
            O => \N__20468\,
            I => \il_max_comp2_D1\
        );

    \I__2465\ : InMux
    port map (
            O => \N__20465\,
            I => \N__20462\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__20462\,
            I => \N__20459\
        );

    \I__2463\ : Glb2LocalMux
    port map (
            O => \N__20459\,
            I => \N__20456\
        );

    \I__2462\ : GlobalMux
    port map (
            O => \N__20456\,
            I => clk_12mhz
        );

    \I__2461\ : IoInMux
    port map (
            O => \N__20453\,
            I => \N__20450\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__20450\,
            I => \N__20447\
        );

    \I__2459\ : IoSpan4Mux
    port map (
            O => \N__20447\,
            I => \N__20444\
        );

    \I__2458\ : Span4Mux_s0_v
    port map (
            O => \N__20444\,
            I => \N__20441\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__20441\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2456\ : InMux
    port map (
            O => \N__20438\,
            I => \N__20435\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__20435\,
            I => \N__20432\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__20432\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__2452\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20423\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__20423\,
            I => \N__20420\
        );

    \I__2450\ : Span4Mux_h
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__20417\,
            I => \current_shift_inst.PI_CTRL.N_155\
        );

    \I__2448\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__20408\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2445\ : InMux
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__20402\,
            I => \N__20399\
        );

    \I__2443\ : Odrv12
    port map (
            O => \N__20399\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2442\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__20390\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9\
        );

    \I__2439\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20384\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__20381\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__2436\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20373\
        );

    \I__2435\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20370\
        );

    \I__2434\ : InMux
    port map (
            O => \N__20376\,
            I => \N__20367\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__20373\,
            I => \N__20364\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__20370\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__20367\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__20364\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__20357\,
            I => \N__20354\
        );

    \I__2428\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__20351\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2426\ : InMux
    port map (
            O => \N__20348\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2425\ : IoInMux
    port map (
            O => \N__20345\,
            I => \N__20342\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__2423\ : IoSpan4Mux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__2422\ : Sp12to4
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__2421\ : Span12Mux_s9_v
    port map (
            O => \N__20333\,
            I => \N__20330\
        );

    \I__2420\ : Span12Mux_h
    port map (
            O => \N__20330\,
            I => \N__20327\
        );

    \I__2419\ : Odrv12
    port map (
            O => \N__20327\,
            I => pwm_output_c
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__20324\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__20321\,
            I => \N__20316\
        );

    \I__2416\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20312\
        );

    \I__2415\ : InMux
    port map (
            O => \N__20319\,
            I => \N__20305\
        );

    \I__2414\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20305\
        );

    \I__2413\ : InMux
    port map (
            O => \N__20315\,
            I => \N__20302\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__20312\,
            I => \N__20299\
        );

    \I__2411\ : InMux
    port map (
            O => \N__20311\,
            I => \N__20294\
        );

    \I__2410\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20294\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__20305\,
            I => \N__20291\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__20302\,
            I => \N__20287\
        );

    \I__2407\ : Span4Mux_h
    port map (
            O => \N__20299\,
            I => \N__20284\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__20294\,
            I => \N__20279\
        );

    \I__2405\ : Span4Mux_h
    port map (
            O => \N__20291\,
            I => \N__20279\
        );

    \I__2404\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20276\
        );

    \I__2403\ : Odrv12
    port map (
            O => \N__20287\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__20284\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__20279\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__20276\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2399\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20264\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__20264\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2397\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20258\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__20258\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__20255\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\
        );

    \I__2394\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20249\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__20249\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__2392\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20242\
        );

    \I__2391\ : InMux
    port map (
            O => \N__20245\,
            I => \N__20238\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__20242\,
            I => \N__20235\
        );

    \I__2389\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20232\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__20238\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2387\ : Odrv4
    port map (
            O => \N__20235\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__20232\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__20225\,
            I => \N__20222\
        );

    \I__2384\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__20219\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2382\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20213\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__20213\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__2380\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20205\
        );

    \I__2379\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20202\
        );

    \I__2378\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20199\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__20205\,
            I => \N__20196\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__20202\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__20199\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__20196\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__20189\,
            I => \N__20186\
        );

    \I__2372\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__20183\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2370\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20176\
        );

    \I__2369\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20172\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__20176\,
            I => \N__20169\
        );

    \I__2367\ : InMux
    port map (
            O => \N__20175\,
            I => \N__20166\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__20172\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__20169\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__20166\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2363\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20156\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__20156\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__20153\,
            I => \N__20150\
        );

    \I__2360\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20147\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__20147\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2358\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20141\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__20141\,
            I => \N__20138\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__20138\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__2355\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20131\
        );

    \I__2354\ : InMux
    port map (
            O => \N__20134\,
            I => \N__20127\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__20131\,
            I => \N__20124\
        );

    \I__2352\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20121\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__20127\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__20124\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__20121\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__2347\ : InMux
    port map (
            O => \N__20111\,
            I => \N__20108\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__20108\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2345\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__20102\,
            I => \N__20097\
        );

    \I__2343\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20094\
        );

    \I__2342\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20091\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__20097\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__20094\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__20091\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2338\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__20081\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__2335\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20072\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__20072\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2333\ : InMux
    port map (
            O => \N__20069\,
            I => \N__20066\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__2331\ : Span4Mux_h
    port map (
            O => \N__20063\,
            I => \N__20060\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__20060\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__2329\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20054\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__20054\,
            I => \N__20049\
        );

    \I__2327\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20046\
        );

    \I__2326\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20043\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__20049\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__20046\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__20043\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__2321\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__20030\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2319\ : InMux
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__2317\ : Odrv12
    port map (
            O => \N__20021\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__2316\ : InMux
    port map (
            O => \N__20018\,
            I => \N__20014\
        );

    \I__2315\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20010\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__20007\
        );

    \I__2313\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20004\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__20010\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__20007\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__20004\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2309\ : CascadeMux
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__2308\ : InMux
    port map (
            O => \N__19994\,
            I => \N__19991\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__19991\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2306\ : InMux
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__2304\ : Odrv12
    port map (
            O => \N__19982\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__2303\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19974\
        );

    \I__2302\ : InMux
    port map (
            O => \N__19978\,
            I => \N__19971\
        );

    \I__2301\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19968\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__19974\,
            I => \N__19965\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__19971\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__19968\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__19965\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__2295\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19952\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__19952\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__19949\,
            I => \N__19946\
        );

    \I__2292\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19941\
        );

    \I__2291\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19936\
        );

    \I__2290\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19936\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__19941\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__19936\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2287\ : InMux
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__2285\ : Odrv12
    port map (
            O => \N__19925\,
            I => il_max_comp2_c
        );

    \I__2284\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__19916\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__2281\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19910\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__19910\,
            I => \N__19907\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__19907\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__2278\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__2276\ : Odrv12
    port map (
            O => \N__19898\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__2275\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__19889\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__2272\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__19883\,
            I => \N__19880\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__19880\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__2268\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__19871\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__2266\ : InMux
    port map (
            O => \N__19868\,
            I => \N__19863\
        );

    \I__2265\ : InMux
    port map (
            O => \N__19867\,
            I => \N__19860\
        );

    \I__2264\ : InMux
    port map (
            O => \N__19866\,
            I => \N__19857\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__19863\,
            I => \N__19854\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__19860\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__19857\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__19854\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2259\ : InMux
    port map (
            O => \N__19847\,
            I => \N__19844\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__19844\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__19841\,
            I => \N__19837\
        );

    \I__2256\ : InMux
    port map (
            O => \N__19840\,
            I => \N__19834\
        );

    \I__2255\ : InMux
    port map (
            O => \N__19837\,
            I => \N__19831\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__19834\,
            I => \N__19828\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__19831\,
            I => \N__19823\
        );

    \I__2252\ : Span4Mux_v
    port map (
            O => \N__19828\,
            I => \N__19823\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__19823\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__2250\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__19817\,
            I => \N__19813\
        );

    \I__2248\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19809\
        );

    \I__2247\ : Span4Mux_h
    port map (
            O => \N__19813\,
            I => \N__19806\
        );

    \I__2246\ : InMux
    port map (
            O => \N__19812\,
            I => \N__19803\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__19809\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__19806\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__19803\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__19796\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\
        );

    \I__2241\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__19790\,
            I => \N__19786\
        );

    \I__2239\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19783\
        );

    \I__2238\ : Span4Mux_v
    port map (
            O => \N__19786\,
            I => \N__19777\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__19783\,
            I => \N__19777\
        );

    \I__2236\ : InMux
    port map (
            O => \N__19782\,
            I => \N__19774\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__19777\,
            I => pwm_duty_input_9
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__19774\,
            I => pwm_duty_input_9
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__19769\,
            I => \N__19764\
        );

    \I__2232\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19761\
        );

    \I__2231\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19758\
        );

    \I__2230\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19755\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__19761\,
            I => \N__19752\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__19758\,
            I => \N__19749\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__19755\,
            I => \N__19742\
        );

    \I__2226\ : Span4Mux_v
    port map (
            O => \N__19752\,
            I => \N__19742\
        );

    \I__2225\ : Span4Mux_v
    port map (
            O => \N__19749\,
            I => \N__19742\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__19742\,
            I => pwm_duty_input_6
        );

    \I__2223\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19734\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__19738\,
            I => \N__19731\
        );

    \I__2221\ : InMux
    port map (
            O => \N__19737\,
            I => \N__19728\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__19734\,
            I => \N__19725\
        );

    \I__2219\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19722\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__19728\,
            I => \N__19719\
        );

    \I__2217\ : Span4Mux_h
    port map (
            O => \N__19725\,
            I => \N__19716\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__19722\,
            I => \N__19711\
        );

    \I__2215\ : Span4Mux_h
    port map (
            O => \N__19719\,
            I => \N__19711\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__19716\,
            I => pwm_duty_input_7
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__19711\,
            I => pwm_duty_input_7
        );

    \I__2212\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19702\
        );

    \I__2211\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19699\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__19702\,
            I => \N__19696\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__19699\,
            I => \N__19693\
        );

    \I__2208\ : Span4Mux_h
    port map (
            O => \N__19696\,
            I => \N__19689\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__19693\,
            I => \N__19686\
        );

    \I__2206\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19683\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__19689\,
            I => pwm_duty_input_8
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__19686\,
            I => pwm_duty_input_8
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__19683\,
            I => pwm_duty_input_8
        );

    \I__2202\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__19670\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\
        );

    \I__2199\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__2197\ : Odrv4
    port map (
            O => \N__19661\,
            I => \current_shift_inst.PI_CTRL.N_149\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__2195\ : InMux
    port map (
            O => \N__19655\,
            I => \N__19651\
        );

    \I__2194\ : InMux
    port map (
            O => \N__19654\,
            I => \N__19648\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__19651\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__19648\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2191\ : CascadeMux
    port map (
            O => \N__19643\,
            I => \N__19637\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__19642\,
            I => \N__19634\
        );

    \I__2189\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19624\
        );

    \I__2188\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19624\
        );

    \I__2187\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19624\
        );

    \I__2186\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19624\
        );

    \I__2185\ : InMux
    port map (
            O => \N__19633\,
            I => \N__19621\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__19624\,
            I => \N__19618\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19615\
        );

    \I__2182\ : Odrv12
    port map (
            O => \N__19618\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__19615\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__19610\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__2179\ : InMux
    port map (
            O => \N__19607\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__2178\ : InMux
    port map (
            O => \N__19604\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__2177\ : InMux
    port map (
            O => \N__19601\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__2176\ : InMux
    port map (
            O => \N__19598\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__2175\ : InMux
    port map (
            O => \N__19595\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__2174\ : InMux
    port map (
            O => \N__19592\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__2173\ : InMux
    port map (
            O => \N__19589\,
            I => \bfn_4_10_0_\
        );

    \I__2172\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19568\
        );

    \I__2171\ : InMux
    port map (
            O => \N__19585\,
            I => \N__19568\
        );

    \I__2170\ : InMux
    port map (
            O => \N__19584\,
            I => \N__19568\
        );

    \I__2169\ : InMux
    port map (
            O => \N__19583\,
            I => \N__19568\
        );

    \I__2168\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19563\
        );

    \I__2167\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19563\
        );

    \I__2166\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19554\
        );

    \I__2165\ : InMux
    port map (
            O => \N__19579\,
            I => \N__19554\
        );

    \I__2164\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19554\
        );

    \I__2163\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19554\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__19568\,
            I => \N__19547\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__19563\,
            I => \N__19547\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__19554\,
            I => \N__19547\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__19547\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2158\ : InMux
    port map (
            O => \N__19544\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__2157\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19537\
        );

    \I__2156\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19534\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__19537\,
            I => \N__19531\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__19534\,
            I => \N__19527\
        );

    \I__2153\ : Span4Mux_v
    port map (
            O => \N__19531\,
            I => \N__19524\
        );

    \I__2152\ : InMux
    port map (
            O => \N__19530\,
            I => \N__19521\
        );

    \I__2151\ : Span4Mux_h
    port map (
            O => \N__19527\,
            I => \N__19518\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__19524\,
            I => pwm_duty_input_4
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__19521\,
            I => pwm_duty_input_4
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__19518\,
            I => pwm_duty_input_4
        );

    \I__2147\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__19505\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__2144\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19488\
        );

    \I__2143\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19488\
        );

    \I__2142\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19483\
        );

    \I__2141\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19483\
        );

    \I__2140\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19480\
        );

    \I__2139\ : InMux
    port map (
            O => \N__19497\,
            I => \N__19469\
        );

    \I__2138\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19469\
        );

    \I__2137\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19469\
        );

    \I__2136\ : InMux
    port map (
            O => \N__19494\,
            I => \N__19469\
        );

    \I__2135\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19469\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__19488\,
            I => \N__19466\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__19483\,
            I => \N__19463\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__19480\,
            I => \N__19460\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__19469\,
            I => \N__19457\
        );

    \I__2130\ : Span4Mux_s3_h
    port map (
            O => \N__19466\,
            I => \N__19450\
        );

    \I__2129\ : Span4Mux_v
    port map (
            O => \N__19463\,
            I => \N__19450\
        );

    \I__2128\ : Span4Mux_h
    port map (
            O => \N__19460\,
            I => \N__19450\
        );

    \I__2127\ : Odrv12
    port map (
            O => \N__19457\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__19450\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__19445\,
            I => \N__19437\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__19444\,
            I => \N__19434\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__19443\,
            I => \N__19428\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__19442\,
            I => \N__19425\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__19441\,
            I => \N__19422\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__19440\,
            I => \N__19419\
        );

    \I__2119\ : InMux
    port map (
            O => \N__19437\,
            I => \N__19406\
        );

    \I__2118\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19406\
        );

    \I__2117\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19403\
        );

    \I__2116\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19392\
        );

    \I__2115\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19392\
        );

    \I__2114\ : InMux
    port map (
            O => \N__19428\,
            I => \N__19392\
        );

    \I__2113\ : InMux
    port map (
            O => \N__19425\,
            I => \N__19392\
        );

    \I__2112\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19392\
        );

    \I__2111\ : InMux
    port map (
            O => \N__19419\,
            I => \N__19387\
        );

    \I__2110\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19387\
        );

    \I__2109\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19382\
        );

    \I__2108\ : InMux
    port map (
            O => \N__19416\,
            I => \N__19382\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__19415\,
            I => \N__19379\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__19414\,
            I => \N__19376\
        );

    \I__2105\ : InMux
    port map (
            O => \N__19413\,
            I => \N__19369\
        );

    \I__2104\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19369\
        );

    \I__2103\ : InMux
    port map (
            O => \N__19411\,
            I => \N__19369\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__19406\,
            I => \N__19366\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__19403\,
            I => \N__19346\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__19392\,
            I => \N__19346\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__19387\,
            I => \N__19341\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__19382\,
            I => \N__19341\
        );

    \I__2097\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19336\
        );

    \I__2096\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19336\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__19369\,
            I => \N__19333\
        );

    \I__2094\ : Span4Mux_h
    port map (
            O => \N__19366\,
            I => \N__19330\
        );

    \I__2093\ : InMux
    port map (
            O => \N__19365\,
            I => \N__19313\
        );

    \I__2092\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19313\
        );

    \I__2091\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19313\
        );

    \I__2090\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19313\
        );

    \I__2089\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19313\
        );

    \I__2088\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19313\
        );

    \I__2087\ : InMux
    port map (
            O => \N__19359\,
            I => \N__19313\
        );

    \I__2086\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19313\
        );

    \I__2085\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19298\
        );

    \I__2084\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19298\
        );

    \I__2083\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19298\
        );

    \I__2082\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19298\
        );

    \I__2081\ : InMux
    port map (
            O => \N__19353\,
            I => \N__19298\
        );

    \I__2080\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19298\
        );

    \I__2079\ : InMux
    port map (
            O => \N__19351\,
            I => \N__19298\
        );

    \I__2078\ : Span4Mux_h
    port map (
            O => \N__19346\,
            I => \N__19293\
        );

    \I__2077\ : Span4Mux_v
    port map (
            O => \N__19341\,
            I => \N__19293\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__19336\,
            I => \N__19288\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__19333\,
            I => \N__19288\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__19330\,
            I => \N_19_1\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__19313\,
            I => \N_19_1\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__19298\,
            I => \N_19_1\
        );

    \I__2071\ : Odrv4
    port map (
            O => \N__19293\,
            I => \N_19_1\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__19288\,
            I => \N_19_1\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__2068\ : InMux
    port map (
            O => \N__19274\,
            I => \N__19271\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__19268\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__2065\ : InMux
    port map (
            O => \N__19265\,
            I => \N__19259\
        );

    \I__2064\ : InMux
    port map (
            O => \N__19264\,
            I => \N__19259\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__19259\,
            I => \N__19250\
        );

    \I__2062\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19247\
        );

    \I__2061\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19236\
        );

    \I__2060\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19236\
        );

    \I__2059\ : InMux
    port map (
            O => \N__19255\,
            I => \N__19236\
        );

    \I__2058\ : InMux
    port map (
            O => \N__19254\,
            I => \N__19236\
        );

    \I__2057\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19236\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__19250\,
            I => \N__19227\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__19247\,
            I => \N__19227\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__19236\,
            I => \N__19227\
        );

    \I__2053\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19222\
        );

    \I__2052\ : InMux
    port map (
            O => \N__19234\,
            I => \N__19222\
        );

    \I__2051\ : Span4Mux_v
    port map (
            O => \N__19227\,
            I => \N__19219\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__19222\,
            I => \N__19216\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__19219\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2048\ : Odrv12
    port map (
            O => \N__19216\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2047\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__19208\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__2045\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__19199\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__2042\ : InMux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__19193\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__2040\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__19187\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__2038\ : InMux
    port map (
            O => \N__19184\,
            I => \bfn_4_9_0_\
        );

    \I__2037\ : InMux
    port map (
            O => \N__19181\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__2036\ : InMux
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__19175\,
            I => \N__19171\
        );

    \I__2034\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19168\
        );

    \I__2033\ : Span4Mux_h
    port map (
            O => \N__19171\,
            I => \N__19165\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__19168\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__19165\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__2030\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__19157\,
            I => \N__19152\
        );

    \I__2028\ : InMux
    port map (
            O => \N__19156\,
            I => \N__19149\
        );

    \I__2027\ : InMux
    port map (
            O => \N__19155\,
            I => \N__19146\
        );

    \I__2026\ : Span4Mux_s3_h
    port map (
            O => \N__19152\,
            I => \N__19141\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__19149\,
            I => \N__19141\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__19146\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__19141\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2022\ : InMux
    port map (
            O => \N__19136\,
            I => \N__19133\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__19133\,
            I => \N__19129\
        );

    \I__2020\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19126\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__19129\,
            I => pwm_duty_input_0
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__19126\,
            I => pwm_duty_input_0
        );

    \I__2017\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__19118\,
            I => \N__19114\
        );

    \I__2015\ : InMux
    port map (
            O => \N__19117\,
            I => \N__19111\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__19114\,
            I => pwm_duty_input_1
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__19111\,
            I => pwm_duty_input_1
        );

    \I__2012\ : InMux
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__19103\,
            I => \N__19099\
        );

    \I__2010\ : InMux
    port map (
            O => \N__19102\,
            I => \N__19096\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__19099\,
            I => pwm_duty_input_2
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__19096\,
            I => pwm_duty_input_2
        );

    \I__2007\ : InMux
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__19088\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__2005\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19081\
        );

    \I__2004\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19078\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__19081\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__19078\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2001\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19067\
        );

    \I__2000\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19067\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__1998\ : Span4Mux_h
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__19061\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1996\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19055\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__19055\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__19052\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__19049\,
            I => \N__19042\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__19048\,
            I => \N__19039\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__19047\,
            I => \N__19036\
        );

    \I__1990\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19033\
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__19045\,
            I => \N__19030\
        );

    \I__1988\ : InMux
    port map (
            O => \N__19042\,
            I => \N__19023\
        );

    \I__1987\ : InMux
    port map (
            O => \N__19039\,
            I => \N__19023\
        );

    \I__1986\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19019\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__19033\,
            I => \N__19015\
        );

    \I__1984\ : InMux
    port map (
            O => \N__19030\,
            I => \N__19008\
        );

    \I__1983\ : InMux
    port map (
            O => \N__19029\,
            I => \N__19008\
        );

    \I__1982\ : InMux
    port map (
            O => \N__19028\,
            I => \N__19008\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__19023\,
            I => \N__19003\
        );

    \I__1980\ : InMux
    port map (
            O => \N__19022\,
            I => \N__19000\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__19019\,
            I => \N__18997\
        );

    \I__1978\ : InMux
    port map (
            O => \N__19018\,
            I => \N__18994\
        );

    \I__1977\ : Span4Mux_h
    port map (
            O => \N__19015\,
            I => \N__18989\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__19008\,
            I => \N__18989\
        );

    \I__1975\ : InMux
    port map (
            O => \N__19007\,
            I => \N__18984\
        );

    \I__1974\ : InMux
    port map (
            O => \N__19006\,
            I => \N__18984\
        );

    \I__1973\ : Span4Mux_s3_h
    port map (
            O => \N__19003\,
            I => \N__18979\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__19000\,
            I => \N__18979\
        );

    \I__1971\ : Odrv12
    port map (
            O => \N__18997\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__18994\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__18989\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__18984\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__18979\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__1966\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18965\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__18965\,
            I => \N__18962\
        );

    \I__1964\ : Span4Mux_v
    port map (
            O => \N__18962\,
            I => \N__18959\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__18959\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__1962\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18953\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__18953\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__18950\,
            I => \N__18947\
        );

    \I__1959\ : InMux
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__18944\,
            I => \N__18941\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__18941\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__18938\,
            I => \N__18935\
        );

    \I__1955\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18931\
        );

    \I__1954\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18928\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__18931\,
            I => \N__18925\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__18928\,
            I => \N__18922\
        );

    \I__1951\ : Span4Mux_h
    port map (
            O => \N__18925\,
            I => \N__18919\
        );

    \I__1950\ : Span4Mux_h
    port map (
            O => \N__18922\,
            I => \N__18916\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__18919\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__18916\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1947\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18906\
        );

    \I__1946\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18903\
        );

    \I__1945\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18900\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__18906\,
            I => \N__18897\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__18903\,
            I => \N__18894\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__18900\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__18897\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1940\ : Odrv12
    port map (
            O => \N__18894\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1939\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__18884\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__1937\ : InMux
    port map (
            O => \N__18881\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__1936\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__18875\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__1934\ : InMux
    port map (
            O => \N__18872\,
            I => \bfn_3_11_0_\
        );

    \I__1933\ : InMux
    port map (
            O => \N__18869\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__1932\ : InMux
    port map (
            O => \N__18866\,
            I => \N__18861\
        );

    \I__1931\ : InMux
    port map (
            O => \N__18865\,
            I => \N__18858\
        );

    \I__1930\ : InMux
    port map (
            O => \N__18864\,
            I => \N__18855\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__18861\,
            I => \N__18852\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__18858\,
            I => \N__18849\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__18855\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__18852\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__18849\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__1924\ : InMux
    port map (
            O => \N__18842\,
            I => \N__18839\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__18839\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__1922\ : InMux
    port map (
            O => \N__18836\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__1921\ : InMux
    port map (
            O => \N__18833\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__1920\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__18824\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__1917\ : InMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__18818\,
            I => \N__18814\
        );

    \I__1915\ : InMux
    port map (
            O => \N__18817\,
            I => \N__18810\
        );

    \I__1914\ : Span4Mux_h
    port map (
            O => \N__18814\,
            I => \N__18807\
        );

    \I__1913\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18804\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__18810\,
            I => pwm_duty_input_3
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__18807\,
            I => pwm_duty_input_3
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__18804\,
            I => pwm_duty_input_3
        );

    \I__1909\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18793\
        );

    \I__1908\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18790\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__18793\,
            I => \N__18787\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__18790\,
            I => \N__18784\
        );

    \I__1905\ : Span4Mux_h
    port map (
            O => \N__18787\,
            I => \N__18781\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__18784\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__18781\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__1901\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18768\
        );

    \I__1900\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18763\
        );

    \I__1899\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18763\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__18768\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__18763\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__1896\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__18755\,
            I => \N__18751\
        );

    \I__1894\ : InMux
    port map (
            O => \N__18754\,
            I => \N__18748\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__18751\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__18748\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1891\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18734\
        );

    \I__1890\ : InMux
    port map (
            O => \N__18742\,
            I => \N__18734\
        );

    \I__1889\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18734\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__18734\,
            I => \N__18731\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__18731\,
            I => \current_shift_inst.PI_CTRL.N_154\
        );

    \I__1886\ : InMux
    port map (
            O => \N__18728\,
            I => \N__18725\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__18725\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \I__1884\ : InMux
    port map (
            O => \N__18722\,
            I => \N__18719\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__18719\,
            I => \N__18716\
        );

    \I__1882\ : Span4Mux_v
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__18713\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1880\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__18707\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__1878\ : InMux
    port map (
            O => \N__18704\,
            I => \N__18701\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__18701\,
            I => \N__18698\
        );

    \I__1876\ : Span4Mux_v
    port map (
            O => \N__18698\,
            I => \N__18695\
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__18695\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1874\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__18689\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__1872\ : InMux
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__18683\,
            I => \N__18680\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__18680\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__1869\ : InMux
    port map (
            O => \N__18677\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__1868\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__18671\,
            I => \N__18667\
        );

    \I__1866\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18664\
        );

    \I__1865\ : Span4Mux_h
    port map (
            O => \N__18667\,
            I => \N__18661\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__18664\,
            I => \N__18658\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__18661\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__18658\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1861\ : InMux
    port map (
            O => \N__18653\,
            I => \N__18650\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__18650\,
            I => \N__18647\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__18647\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__1858\ : InMux
    port map (
            O => \N__18644\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__1857\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18636\
        );

    \I__1856\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18633\
        );

    \I__1855\ : InMux
    port map (
            O => \N__18639\,
            I => \N__18630\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__18636\,
            I => \N__18627\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__18633\,
            I => \N__18624\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__18630\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__18627\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__18624\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1849\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__18614\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__1847\ : InMux
    port map (
            O => \N__18611\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__1846\ : InMux
    port map (
            O => \N__18608\,
            I => \N__18605\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__18605\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__1844\ : InMux
    port map (
            O => \N__18602\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__1843\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__18596\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__1841\ : InMux
    port map (
            O => \N__18593\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__1840\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18583\
        );

    \I__1839\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18583\
        );

    \I__1838\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18580\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__18583\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__18580\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1835\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__18569\,
            I => \N__18566\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__18566\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1831\ : InMux
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__18560\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__1829\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__18548\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1825\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__18542\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__1823\ : InMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__18536\,
            I => \N__18533\
        );

    \I__1821\ : Span4Mux_h
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__18530\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1819\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__18524\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__1817\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__1815\ : Span4Mux_h
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__18512\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1813\ : InMux
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__18506\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__1811\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__1809\ : Span4Mux_h
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__18494\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1807\ : InMux
    port map (
            O => \N__18491\,
            I => \N__18488\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__18488\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__1805\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__1803\ : Span4Mux_h
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__18476\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1801\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__18470\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__1799\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__18464\,
            I => \N__18461\
        );

    \I__1797\ : Span4Mux_h
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__18458\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1795\ : InMux
    port map (
            O => \N__18455\,
            I => \N__18452\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__18452\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__1793\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__1791\ : Span4Mux_h
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__18440\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__18437\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__18434\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__1787\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__18428\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__1785\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__18422\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__1783\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__18416\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__1781\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__18410\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__1778\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__18401\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__1776\ : InMux
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__18395\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__1773\ : InMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__18386\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__1771\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__18380\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__1769\ : CascadeMux
    port map (
            O => \N__18377\,
            I => \N__18368\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__18376\,
            I => \N__18365\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__18375\,
            I => \N__18362\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__18374\,
            I => \N__18358\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__18373\,
            I => \N__18355\
        );

    \I__1764\ : InMux
    port map (
            O => \N__18372\,
            I => \N__18350\
        );

    \I__1763\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18350\
        );

    \I__1762\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18345\
        );

    \I__1761\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18345\
        );

    \I__1760\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18336\
        );

    \I__1759\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18336\
        );

    \I__1758\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18336\
        );

    \I__1757\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18336\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__18350\,
            I => \N__18329\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__18345\,
            I => \N__18329\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__18336\,
            I => \N__18329\
        );

    \I__1753\ : Span4Mux_h
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__18326\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1751\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__18320\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__1749\ : InMux
    port map (
            O => \N__18317\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__1748\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18311\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__18311\,
            I => \N__18308\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__18308\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__1745\ : InMux
    port map (
            O => \N__18305\,
            I => \N__18302\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__18302\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__1743\ : InMux
    port map (
            O => \N__18299\,
            I => \bfn_2_12_0_\
        );

    \I__1742\ : InMux
    port map (
            O => \N__18296\,
            I => \N__18293\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__18293\,
            I => \N__18289\
        );

    \I__1740\ : InMux
    port map (
            O => \N__18292\,
            I => \N__18286\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__18289\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__18286\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__18281\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__18278\,
            I => \N__18275\
        );

    \I__1735\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18272\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__18272\,
            I => \N__18269\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__18269\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__1732\ : InMux
    port map (
            O => \N__18266\,
            I => \N__18257\
        );

    \I__1731\ : InMux
    port map (
            O => \N__18265\,
            I => \N__18257\
        );

    \I__1730\ : InMux
    port map (
            O => \N__18264\,
            I => \N__18257\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__18257\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1728\ : InMux
    port map (
            O => \N__18254\,
            I => \N__18251\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__18251\,
            I => \N__18248\
        );

    \I__1726\ : Odrv12
    port map (
            O => \N__18248\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__1725\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18242\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__18242\,
            I => \N__18239\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__18239\,
            I => \N__18236\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__18236\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__18233\,
            I => \N__18228\
        );

    \I__1720\ : InMux
    port map (
            O => \N__18232\,
            I => \N__18225\
        );

    \I__1719\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18222\
        );

    \I__1718\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18219\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__18225\,
            I => \N__18216\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__18222\,
            I => \N__18213\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__18219\,
            I => \N__18210\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__18216\,
            I => \N__18207\
        );

    \I__1713\ : Span4Mux_v
    port map (
            O => \N__18213\,
            I => \N__18204\
        );

    \I__1712\ : Odrv12
    port map (
            O => \N__18210\,
            I => pwm_duty_input_5
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__18207\,
            I => pwm_duty_input_5
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__18204\,
            I => pwm_duty_input_5
        );

    \I__1709\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18194\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__18194\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__1707\ : InMux
    port map (
            O => \N__18191\,
            I => \N__18188\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__1705\ : Span4Mux_h
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__1704\ : Span4Mux_v
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__18179\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__1701\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__18170\,
            I => \N__18167\
        );

    \I__1699\ : Span4Mux_h
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__18164\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__1697\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__18158\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__1695\ : InMux
    port map (
            O => \N__18155\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__1694\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__18149\,
            I => \N__18146\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__18146\,
            I => \N__18143\
        );

    \I__1691\ : Span4Mux_v
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__18140\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__18137\,
            I => \N__18134\
        );

    \I__1688\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18131\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__18131\,
            I => \N__18128\
        );

    \I__1686\ : Span4Mux_h
    port map (
            O => \N__18128\,
            I => \N__18125\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__18125\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__1684\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18119\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__18119\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__1682\ : InMux
    port map (
            O => \N__18116\,
            I => \bfn_2_11_0_\
        );

    \I__1681\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18110\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__18110\,
            I => \N__18107\
        );

    \I__1679\ : Span4Mux_h
    port map (
            O => \N__18107\,
            I => \N__18104\
        );

    \I__1678\ : Span4Mux_v
    port map (
            O => \N__18104\,
            I => \N__18101\
        );

    \I__1677\ : Odrv4
    port map (
            O => \N__18101\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__18098\,
            I => \N__18095\
        );

    \I__1675\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__18092\,
            I => \N__18089\
        );

    \I__1673\ : Span4Mux_h
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__1672\ : Span4Mux_s0_h
    port map (
            O => \N__18086\,
            I => \N__18083\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__18083\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__1670\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18077\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__18077\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__1668\ : InMux
    port map (
            O => \N__18074\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1667\ : InMux
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__1665\ : Span4Mux_h
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__1664\ : Span4Mux_v
    port map (
            O => \N__18062\,
            I => \N__18059\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__18059\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1662\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__18053\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__1660\ : InMux
    port map (
            O => \N__18050\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1659\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18044\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__18038\,
            I => \N__18035\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__18035\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1654\ : InMux
    port map (
            O => \N__18032\,
            I => \N__18029\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__18029\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__1652\ : InMux
    port map (
            O => \N__18026\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1651\ : InMux
    port map (
            O => \N__18023\,
            I => \N__18020\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__18020\,
            I => \N__18017\
        );

    \I__1649\ : Span4Mux_v
    port map (
            O => \N__18017\,
            I => \N__18014\
        );

    \I__1648\ : Span4Mux_v
    port map (
            O => \N__18014\,
            I => \N__18011\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__18011\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1646\ : InMux
    port map (
            O => \N__18008\,
            I => \N__18005\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__18005\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__1644\ : InMux
    port map (
            O => \N__18002\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__1642\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17993\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__17993\,
            I => \N__17990\
        );

    \I__1640\ : Span12Mux_h
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__1639\ : Odrv12
    port map (
            O => \N__17987\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__1638\ : InMux
    port map (
            O => \N__17984\,
            I => \N__17981\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__17981\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__1636\ : InMux
    port map (
            O => \N__17978\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__1635\ : InMux
    port map (
            O => \N__17975\,
            I => \N__17972\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__17972\,
            I => \N__17969\
        );

    \I__1633\ : Span12Mux_v
    port map (
            O => \N__17969\,
            I => \N__17966\
        );

    \I__1632\ : Odrv12
    port map (
            O => \N__17966\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__1631\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17960\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__17960\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__1629\ : InMux
    port map (
            O => \N__17957\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__1628\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17951\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__17951\,
            I => \N__17948\
        );

    \I__1626\ : Span4Mux_h
    port map (
            O => \N__17948\,
            I => \N__17945\
        );

    \I__1625\ : Span4Mux_v
    port map (
            O => \N__17945\,
            I => \N__17942\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__17942\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__17939\,
            I => \N__17936\
        );

    \I__1622\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17933\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__17933\,
            I => \N__17930\
        );

    \I__1620\ : Span4Mux_h
    port map (
            O => \N__17930\,
            I => \N__17927\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__17927\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1618\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17921\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__17921\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__1616\ : InMux
    port map (
            O => \N__17918\,
            I => \N__17915\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__17915\,
            I => \N__17912\
        );

    \I__1614\ : Span4Mux_h
    port map (
            O => \N__17912\,
            I => \N__17909\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__17909\,
            I => \N__17906\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__17906\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__17903\,
            I => \N__17900\
        );

    \I__1610\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__17897\,
            I => \N__17894\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__17894\,
            I => \N__17891\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__17891\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__17888\,
            I => \N__17885\
        );

    \I__1605\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17882\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__17882\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__1603\ : InMux
    port map (
            O => \N__17879\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1602\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17873\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__17873\,
            I => \N__17870\
        );

    \I__1600\ : Span4Mux_h
    port map (
            O => \N__17870\,
            I => \N__17867\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__17867\,
            I => \N__17864\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__17864\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__17861\,
            I => \N__17858\
        );

    \I__1596\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17855\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__17855\,
            I => \N__17852\
        );

    \I__1594\ : Span4Mux_h
    port map (
            O => \N__17852\,
            I => \N__17849\
        );

    \I__1593\ : Odrv4
    port map (
            O => \N__17849\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1592\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__17843\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__1590\ : InMux
    port map (
            O => \N__17840\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1589\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__17834\,
            I => \N__17831\
        );

    \I__1587\ : Span4Mux_h
    port map (
            O => \N__17831\,
            I => \N__17828\
        );

    \I__1586\ : Span4Mux_v
    port map (
            O => \N__17828\,
            I => \N__17825\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__17825\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__17822\,
            I => \N__17819\
        );

    \I__1583\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17816\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__17816\,
            I => \N__17813\
        );

    \I__1581\ : Span4Mux_v
    port map (
            O => \N__17813\,
            I => \N__17810\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__17810\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__17807\,
            I => \N__17804\
        );

    \I__1578\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17801\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__17801\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__1576\ : InMux
    port map (
            O => \N__17798\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1575\ : InMux
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__17789\,
            I => \N__17786\
        );

    \I__1572\ : Span4Mux_v
    port map (
            O => \N__17786\,
            I => \N__17783\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__17783\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__17780\,
            I => \N__17777\
        );

    \I__1569\ : InMux
    port map (
            O => \N__17777\,
            I => \N__17774\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__17774\,
            I => \N__17771\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__17771\,
            I => \N__17768\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__17768\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1565\ : InMux
    port map (
            O => \N__17765\,
            I => \N__17762\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__17762\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__1563\ : InMux
    port map (
            O => \N__17759\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1562\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17753\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__17753\,
            I => \N__17750\
        );

    \I__1560\ : Span12Mux_h
    port map (
            O => \N__17750\,
            I => \N__17747\
        );

    \I__1559\ : Odrv12
    port map (
            O => \N__17747\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__17744\,
            I => \N__17741\
        );

    \I__1557\ : InMux
    port map (
            O => \N__17741\,
            I => \N__17738\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__17738\,
            I => \N__17735\
        );

    \I__1555\ : Span4Mux_h
    port map (
            O => \N__17735\,
            I => \N__17732\
        );

    \I__1554\ : Span4Mux_s0_h
    port map (
            O => \N__17732\,
            I => \N__17729\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__17729\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__1552\ : InMux
    port map (
            O => \N__17726\,
            I => \N__17723\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__17723\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__1550\ : InMux
    port map (
            O => \N__17720\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__1549\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__17714\,
            I => \N__17711\
        );

    \I__1547\ : Span12Mux_v
    port map (
            O => \N__17711\,
            I => \N__17708\
        );

    \I__1546\ : Odrv12
    port map (
            O => \N__17708\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__17705\,
            I => \N__17702\
        );

    \I__1544\ : InMux
    port map (
            O => \N__17702\,
            I => \N__17699\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__17699\,
            I => \N__17696\
        );

    \I__1542\ : Span4Mux_h
    port map (
            O => \N__17696\,
            I => \N__17693\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__17693\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__1540\ : InMux
    port map (
            O => \N__17690\,
            I => \N__17687\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__17687\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__1538\ : InMux
    port map (
            O => \N__17684\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__1537\ : InMux
    port map (
            O => \N__17681\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__1536\ : InMux
    port map (
            O => \N__17678\,
            I => \N__17675\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__17675\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__1534\ : InMux
    port map (
            O => \N__17672\,
            I => \bfn_2_9_0_\
        );

    \I__1533\ : InMux
    port map (
            O => \N__17669\,
            I => \N__17666\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__17666\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__1531\ : InMux
    port map (
            O => \N__17663\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__1530\ : InMux
    port map (
            O => \N__17660\,
            I => \N__17657\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__17657\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__1528\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17648\
        );

    \I__1527\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17648\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__17648\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__17645\,
            I => \N__17642\
        );

    \I__1524\ : InMux
    port map (
            O => \N__17642\,
            I => \N__17639\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__17639\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__1522\ : CascadeMux
    port map (
            O => \N__17636\,
            I => \N__17632\
        );

    \I__1521\ : InMux
    port map (
            O => \N__17635\,
            I => \N__17629\
        );

    \I__1520\ : InMux
    port map (
            O => \N__17632\,
            I => \N__17626\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__17629\,
            I => \N__17623\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__17626\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__17623\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1516\ : InMux
    port map (
            O => \N__17618\,
            I => \N__17615\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__17615\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__1514\ : InMux
    port map (
            O => \N__17612\,
            I => \N__17609\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__17609\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__1512\ : InMux
    port map (
            O => \N__17606\,
            I => \N__17603\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__17603\,
            I => \rgb_drv_RNOZ0\
        );

    \I__1510\ : InMux
    port map (
            O => \N__17600\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__1509\ : InMux
    port map (
            O => \N__17597\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__1508\ : InMux
    port map (
            O => \N__17594\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__1507\ : InMux
    port map (
            O => \N__17591\,
            I => \N__17588\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__17588\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__1505\ : InMux
    port map (
            O => \N__17585\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__1504\ : InMux
    port map (
            O => \N__17582\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__1503\ : InMux
    port map (
            O => \N__17579\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__1502\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__17567\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \I__1498\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17560\
        );

    \I__1497\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17557\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__17560\,
            I => \N__17552\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__17557\,
            I => \N__17552\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__17552\,
            I => \N__17549\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__17549\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1492\ : InMux
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__17543\,
            I => \N_38_i_i\
        );

    \I__1490\ : InMux
    port map (
            O => \N__17540\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__1489\ : InMux
    port map (
            O => \N__17537\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__1488\ : InMux
    port map (
            O => \N__17534\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__1487\ : InMux
    port map (
            O => \N__17531\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__1486\ : InMux
    port map (
            O => \N__17528\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__1485\ : InMux
    port map (
            O => \N__17525\,
            I => \bfn_1_10_0_\
        );

    \I__1484\ : InMux
    port map (
            O => \N__17522\,
            I => \N__17519\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__17519\,
            I => \N__17516\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__17516\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1481\ : InMux
    port map (
            O => \N__17513\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__17510\,
            I => \N__17507\
        );

    \I__1479\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17504\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__17504\,
            I => \N__17501\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__17501\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1476\ : InMux
    port map (
            O => \N__17498\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__1475\ : InMux
    port map (
            O => \N__17495\,
            I => \N__17492\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__17492\,
            I => \N__17489\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__17489\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1472\ : InMux
    port map (
            O => \N__17486\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__1471\ : IoInMux
    port map (
            O => \N__17483\,
            I => \N__17480\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__17480\,
            I => \N__17477\
        );

    \I__1469\ : Span4Mux_s3_v
    port map (
            O => \N__17477\,
            I => \N__17474\
        );

    \I__1468\ : Span4Mux_h
    port map (
            O => \N__17474\,
            I => \N__17471\
        );

    \I__1467\ : Sp12to4
    port map (
            O => \N__17471\,
            I => \N__17468\
        );

    \I__1466\ : Span12Mux_v
    port map (
            O => \N__17468\,
            I => \N__17465\
        );

    \I__1465\ : Span12Mux_v
    port map (
            O => \N__17465\,
            I => \N__17462\
        );

    \I__1464\ : Odrv12
    port map (
            O => \N__17462\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1463\ : IoInMux
    port map (
            O => \N__17459\,
            I => \N__17456\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__17456\,
            I => \N__17453\
        );

    \I__1461\ : IoSpan4Mux
    port map (
            O => \N__17453\,
            I => \N__17450\
        );

    \I__1460\ : IoSpan4Mux
    port map (
            O => \N__17450\,
            I => \N__17447\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__17447\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_6\,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_14\,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_22\,
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_18_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_18_21_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_3_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_3_10_0_\
        );

    \IN_MUX_bfv_3_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_3_11_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_18_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_7_0_\
        );

    \IN_MUX_bfv_18_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_18_8_0_\
        );

    \IN_MUX_bfv_18_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_18_9_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_7_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_18_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_13_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_13_27_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_7\,
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_12_12_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17483\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17459\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__27833\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_166_i_g\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__36653\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_434_i_g\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__23633\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_432_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__40376\,
            CLKHFEN => \N__40378\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__40377\,
            RGB2PWM => \N__17546\,
            RGB1 => rgb_g_wire,
            CURREN => \N__40485\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__17606\,
            RGB0PWM => \N__44337\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21677\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44951\,
            ce => 'H',
            sr => \N__44170\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__21670\,
            in1 => \N__20555\,
            in2 => \N__21200\,
            in3 => \N__20320\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44950\,
            ce => 'H',
            sr => \N__44183\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__19501\,
            in1 => \N__17591\,
            in2 => \N__19414\,
            in3 => \N__19234\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44950\,
            ce => 'H',
            sr => \N__44183\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__19502\,
            in1 => \N__17678\,
            in2 => \N__19415\,
            in3 => \N__19235\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44950\,
            ce => 'H',
            sr => \N__44183\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18670\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17522\,
            in2 => \_gnd_net_\,
            in3 => \N__17513\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17510\,
            in3 => \N__17498\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17495\,
            in2 => \_gnd_net_\,
            in3 => \N__17486\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17924\,
            in2 => \_gnd_net_\,
            in3 => \N__17537\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40547\,
            in2 => \N__17888\,
            in3 => \N__17534\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17846\,
            in2 => \N__40607\,
            in3 => \N__17531\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40551\,
            in2 => \N__17807\,
            in3 => \N__17528\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17765\,
            in2 => \_gnd_net_\,
            in3 => \N__17525\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17726\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17690\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18161\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18122\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18080\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18056\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18032\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18008\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17984\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17963\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18323\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17540\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__18372\,
            in1 => \N__17563\,
            in2 => \_gnd_net_\,
            in3 => \N__19418\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__17576\,
            in1 => \N__17564\,
            in2 => \N__19440\,
            in3 => \N__18371\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__19676\,
            in1 => \N__18817\,
            in2 => \N__18233\,
            in3 => \N__19541\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__18741\,
            in1 => \N__18265\,
            in2 => \N__19642\,
            in3 => \N__20963\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44942\,
            ce => 'H',
            sr => \N__44217\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__18742\,
            in1 => \N__18266\,
            in2 => \N__19643\,
            in3 => \N__20948\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44942\,
            ce => 'H',
            sr => \N__44217\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18264\,
            in1 => \N__18743\,
            in2 => \N__20930\,
            in3 => \N__19640\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44942\,
            ce => 'H',
            sr => \N__44217\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__21673\,
            in1 => \N__20547\,
            in2 => \N__21095\,
            in3 => \N__20315\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44942\,
            ce => 'H',
            sr => \N__44217\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__20546\,
            in1 => \N__18758\,
            in2 => \N__21275\,
            in3 => \N__19641\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44942\,
            ce => 'H',
            sr => \N__44217\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__21651\,
            in1 => \N__20554\,
            in2 => \N__21164\,
            in3 => \N__20319\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44939\,
            ce => 'H',
            sr => \N__44224\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100100010"
        )
    port map (
            in0 => \N__20553\,
            in1 => \N__21652\,
            in2 => \N__20321\,
            in3 => \N__21053\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44939\,
            ce => 'H',
            sr => \N__44224\
        );

    \rgb_drv_RNO_0_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__44335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26719\,
            lcout => \N_38_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__44336\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26723\,
            lcout => \rgb_drv_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17635\,
            in2 => \_gnd_net_\,
            in3 => \N__18639\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18245\,
            in2 => \N__19047\,
            in3 => \N__19046\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18653\,
            in2 => \_gnd_net_\,
            in3 => \N__17600\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17618\,
            in2 => \_gnd_net_\,
            in3 => \N__17597\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17645\,
            in3 => \N__17594\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17612\,
            in2 => \_gnd_net_\,
            in3 => \N__17585\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17660\,
            in2 => \_gnd_net_\,
            in3 => \N__17582\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18254\,
            in2 => \_gnd_net_\,
            in3 => \N__17579\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18968\,
            in2 => \_gnd_net_\,
            in3 => \N__17681\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18278\,
            in3 => \N__17672\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__18830\,
            in1 => \N__17669\,
            in2 => \N__19049\,
            in3 => \N__17663\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__17654\,
            in1 => \N__18887\,
            in2 => \N__19045\,
            in3 => \N__18589\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__18590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17653\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__19028\,
            in1 => \N__18608\,
            in2 => \N__19841\,
            in3 => \N__19820\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__18617\,
            in1 => \N__18641\,
            in2 => \N__17636\,
            in3 => \N__19029\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__18864\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18292\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__19160\,
            in1 => \N__18599\,
            in2 => \N__19048\,
            in3 => \N__19174\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17954\,
            in2 => \N__17939\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17918\,
            in2 => \N__17903\,
            in3 => \N__17879\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17876\,
            in2 => \N__17861\,
            in3 => \N__17840\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17837\,
            in2 => \N__17822\,
            in3 => \N__17798\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17795\,
            in2 => \N__17780\,
            in3 => \N__17759\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17756\,
            in2 => \N__17744\,
            in3 => \N__17720\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17717\,
            in2 => \N__17705\,
            in3 => \N__17684\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18191\,
            in2 => \N__18176\,
            in3 => \N__18155\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18152\,
            in2 => \N__18137\,
            in3 => \N__18116\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18113\,
            in2 => \N__18098\,
            in3 => \N__18074\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18071\,
            in2 => \N__18373\,
            in3 => \N__18050\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18047\,
            in2 => \N__18376\,
            in3 => \N__18026\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18023\,
            in2 => \N__18374\,
            in3 => \N__18002\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18361\,
            in2 => \N__17999\,
            in3 => \N__17978\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17975\,
            in2 => \N__18375\,
            in3 => \N__17957\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18383\,
            in2 => \N__18377\,
            in3 => \N__18317\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18314\,
            in1 => \N__18305\,
            in2 => \_gnd_net_\,
            in3 => \N__18299\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__18296\,
            in1 => \N__18865\,
            in2 => \N__18281\,
            in3 => \N__18842\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000010"
        )
    port map (
            in0 => \N__18754\,
            in1 => \N__21274\,
            in2 => \N__20552\,
            in3 => \N__19633\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011110000100"
        )
    port map (
            in0 => \N__18878\,
            in1 => \N__19007\,
            in2 => \N__18776\,
            in3 => \N__18796\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__18686\,
            in1 => \N__18911\,
            in2 => \N__18938\,
            in3 => \N__19006\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19739\,
            in2 => \_gnd_net_\,
            in3 => \N__18232\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__19499\,
            in1 => \N__18197\,
            in2 => \N__19444\,
            in3 => \N__19264\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44949\,
            ce => 'H',
            sr => \N__44162\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20210\,
            in2 => \_gnd_net_\,
            in3 => \N__19868\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__20135\,
            in1 => \N__20180\,
            in2 => \N__18437\,
            in3 => \N__20246\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20057\,
            in1 => \N__20105\,
            in2 => \N__18434\,
            in3 => \N__19511\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__19500\,
            in1 => \N__18431\,
            in2 => \N__19445\,
            in3 => \N__19265\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44949\,
            ce => 'H',
            sr => \N__44162\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__19257\,
            in1 => \N__19497\,
            in2 => \N__19443\,
            in3 => \N__18425\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44947\,
            ce => 'H',
            sr => \N__44171\
        );

    \pwm_generator_inst.threshold_6_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18419\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44947\,
            ce => 'H',
            sr => \N__44171\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__19255\,
            in1 => \N__19496\,
            in2 => \N__19442\,
            in3 => \N__18413\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44947\,
            ce => 'H',
            sr => \N__44171\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__19494\,
            in1 => \N__19432\,
            in2 => \N__18407\,
            in3 => \N__19256\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44947\,
            ce => 'H',
            sr => \N__44171\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__19254\,
            in1 => \N__19495\,
            in2 => \N__19441\,
            in3 => \N__18398\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44947\,
            ce => 'H',
            sr => \N__44171\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__19493\,
            in1 => \N__19431\,
            in2 => \N__18392\,
            in3 => \N__19253\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44947\,
            ce => 'H',
            sr => \N__44171\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18563\,
            in2 => \_gnd_net_\,
            in3 => \N__18575\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18545\,
            in2 => \_gnd_net_\,
            in3 => \N__18557\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18527\,
            in2 => \_gnd_net_\,
            in3 => \N__18539\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18509\,
            in2 => \_gnd_net_\,
            in3 => \N__18521\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18491\,
            in2 => \_gnd_net_\,
            in3 => \N__18503\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18473\,
            in2 => \_gnd_net_\,
            in3 => \N__18485\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18455\,
            in2 => \_gnd_net_\,
            in3 => \N__18467\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18728\,
            in2 => \_gnd_net_\,
            in3 => \N__18449\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18710\,
            in2 => \_gnd_net_\,
            in3 => \N__18722\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_3_10_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18692\,
            in2 => \_gnd_net_\,
            in3 => \N__18704\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18910\,
            in2 => \_gnd_net_\,
            in3 => \N__18677\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__19022\,
            in1 => \N__18674\,
            in2 => \_gnd_net_\,
            in3 => \N__18644\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18640\,
            in2 => \_gnd_net_\,
            in3 => \N__18611\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19812\,
            in2 => \_gnd_net_\,
            in3 => \N__18602\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19156\,
            in2 => \_gnd_net_\,
            in3 => \N__18593\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18588\,
            in2 => \_gnd_net_\,
            in3 => \N__18881\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18771\,
            in2 => \_gnd_net_\,
            in3 => \N__18872\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_3_11_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19084\,
            in2 => \_gnd_net_\,
            in3 => \N__18869\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18866\,
            in2 => \_gnd_net_\,
            in3 => \N__18836\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18833\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__19091\,
            in1 => \N__18821\,
            in2 => \N__18950\,
            in3 => \N__19530\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__18772\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18797\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__19944\,
            in1 => \N__21671\,
            in2 => \_gnd_net_\,
            in3 => \N__21239\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__21672\,
            in1 => \N__19945\,
            in2 => \_gnd_net_\,
            in3 => \N__20534\,
            lcout => \current_shift_inst.PI_CTRL.N_154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19155\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19178\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19136\,
            in1 => \N__19121\,
            in2 => \_gnd_net_\,
            in3 => \N__19106\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19072\,
            in2 => \_gnd_net_\,
            in3 => \N__19085\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__19073\,
            in1 => \N__19058\,
            in2 => \N__19052\,
            in3 => \N__19018\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__19705\,
            in1 => \N__19789\,
            in2 => \N__19769\,
            in3 => \N__18956\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__18909\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18934\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_14_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__24749\,
            in1 => \N__21593\,
            in2 => \N__21938\,
            in3 => \N__26032\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44927\,
            ce => \N__25641\,
            sr => \N__44218\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_19_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__26030\,
            in1 => \N__24480\,
            in2 => \_gnd_net_\,
            in3 => \N__24751\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44927\,
            ce => \N__25641\,
            sr => \N__44218\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_18_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__24748\,
            in1 => \N__26031\,
            in2 => \_gnd_net_\,
            in3 => \N__23381\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44927\,
            ce => \N__25641\,
            sr => \N__44218\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_17_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__26029\,
            in1 => \N__23420\,
            in2 => \_gnd_net_\,
            in3 => \N__24750\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44927\,
            ce => \N__25641\,
            sr => \N__44218\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20378\,
            in1 => \N__19979\,
            in2 => \_gnd_net_\,
            in3 => \N__20018\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_0_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19211\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44945\,
            ce => 'H',
            sr => \N__44163\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__19498\,
            in1 => \N__19433\,
            in2 => \N__19277\,
            in3 => \N__19258\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44945\,
            ce => 'H',
            sr => \N__44163\
        );

    \pwm_generator_inst.threshold_4_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19205\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44945\,
            ce => 'H',
            sr => \N__44163\
        );

    \pwm_generator_inst.threshold_5_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19196\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44945\,
            ce => 'H',
            sr => \N__44163\
        );

    \pwm_generator_inst.threshold_2_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19190\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44945\,
            ce => 'H',
            sr => \N__44163\
        );

    \pwm_generator_inst.counter_0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19577\,
            in1 => \N__19867\,
            in2 => \_gnd_net_\,
            in3 => \N__19184\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__44943\,
            ce => 'H',
            sr => \N__44172\
        );

    \pwm_generator_inst.counter_1_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19583\,
            in1 => \N__20245\,
            in2 => \_gnd_net_\,
            in3 => \N__19181\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__44943\,
            ce => 'H',
            sr => \N__44172\
        );

    \pwm_generator_inst.counter_2_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19578\,
            in1 => \N__20209\,
            in2 => \_gnd_net_\,
            in3 => \N__19607\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__44943\,
            ce => 'H',
            sr => \N__44172\
        );

    \pwm_generator_inst.counter_3_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19584\,
            in1 => \N__20179\,
            in2 => \_gnd_net_\,
            in3 => \N__19604\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__44943\,
            ce => 'H',
            sr => \N__44172\
        );

    \pwm_generator_inst.counter_4_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19579\,
            in1 => \N__20134\,
            in2 => \_gnd_net_\,
            in3 => \N__19601\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__44943\,
            ce => 'H',
            sr => \N__44172\
        );

    \pwm_generator_inst.counter_5_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19585\,
            in1 => \N__20101\,
            in2 => \_gnd_net_\,
            in3 => \N__19598\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__44943\,
            ce => 'H',
            sr => \N__44172\
        );

    \pwm_generator_inst.counter_6_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19580\,
            in1 => \N__20053\,
            in2 => \_gnd_net_\,
            in3 => \N__19595\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__44943\,
            ce => 'H',
            sr => \N__44172\
        );

    \pwm_generator_inst.counter_7_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19586\,
            in1 => \N__20017\,
            in2 => \_gnd_net_\,
            in3 => \N__19592\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__44943\,
            ce => 'H',
            sr => \N__44172\
        );

    \pwm_generator_inst.counter_8_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19582\,
            in1 => \N__19978\,
            in2 => \_gnd_net_\,
            in3 => \N__19589\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__44940\,
            ce => 'H',
            sr => \N__44178\
        );

    \pwm_generator_inst.counter_9_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__20377\,
            in1 => \N__19581\,
            in2 => \_gnd_net_\,
            in3 => \N__19544\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44940\,
            ce => 'H',
            sr => \N__44178\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__19667\,
            in1 => \N__21234\,
            in2 => \N__19658\,
            in3 => \N__20310\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44940\,
            ce => 'H',
            sr => \N__44178\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__20548\,
            in1 => \N__21663\,
            in2 => \N__21128\,
            in3 => \N__20311\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44940\,
            ce => 'H',
            sr => \N__44178\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19840\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21192\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21091\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21126\,
            in1 => \N__21157\,
            in2 => \N__19796\,
            in3 => \N__21048\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19793\,
            in1 => \N__19768\,
            in2 => \N__19738\,
            in3 => \N__19706\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__21238\,
            in1 => \N__21662\,
            in2 => \N__19949\,
            in3 => \N__20525\,
            lcout => \current_shift_inst.PI_CTRL.N_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__21661\,
            in1 => \N__19654\,
            in2 => \N__20429\,
            in3 => \N__20290\,
            lcout => \current_shift_inst.PI_CTRL.N_153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__21193\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21049\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__21127\,
            in1 => \N__21084\,
            in2 => \N__19610\,
            in3 => \N__21150\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19931\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_7_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19922\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44946\,
            ce => 'H',
            sr => \N__44151\
        );

    \pwm_generator_inst.threshold_3_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19913\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44944\,
            ce => 'H',
            sr => \N__44158\
        );

    \pwm_generator_inst.threshold_8_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19904\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44944\,
            ce => 'H',
            sr => \N__44158\
        );

    \pwm_generator_inst.threshold_9_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19895\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44944\,
            ce => 'H',
            sr => \N__44158\
        );

    \pwm_generator_inst.threshold_1_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19886\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44944\,
            ce => 'H',
            sr => \N__44158\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19847\,
            in2 => \N__19877\,
            in3 => \N__19866\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20252\,
            in2 => \N__20225\,
            in3 => \N__20241\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20216\,
            in2 => \N__20189\,
            in3 => \N__20208\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20175\,
            in1 => \N__20159\,
            in2 => \N__20153\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20144\,
            in2 => \N__20114\,
            in3 => \N__20130\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20100\,
            in1 => \N__20084\,
            in2 => \N__20078\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20069\,
            in2 => \N__20036\,
            in3 => \N__20052\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20027\,
            in2 => \N__19997\,
            in3 => \N__20013\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19988\,
            in2 => \N__19958\,
            in3 => \N__19977\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20387\,
            in2 => \N__20357\,
            in3 => \N__20376\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20348\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44936\,
            ce => 'H',
            sr => \N__44173\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20261\,
            in1 => \N__20438\,
            in2 => \N__21416\,
            in3 => \N__21008\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_15_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21482\,
            in1 => \N__21365\,
            in2 => \N__21344\,
            in3 => \N__20396\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20267\,
            in1 => \N__20591\,
            in2 => \N__20324\,
            in3 => \N__20570\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21704\,
            in1 => \N__21461\,
            in2 => \N__21308\,
            in3 => \N__21322\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21304\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20483\,
            in1 => \N__21545\,
            in2 => \N__21566\,
            in3 => \N__21437\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20414\,
            in1 => \N__20405\,
            in2 => \N__20255\,
            in3 => \N__20561\,
            lcout => \current_shift_inst.PI_CTRL.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21700\,
            in2 => \_gnd_net_\,
            in3 => \N__21460\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20477\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44891\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20465\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21409\,
            in2 => \_gnd_net_\,
            in3 => \N__21019\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21020\,
            in1 => \N__21358\,
            in2 => \N__21731\,
            in3 => \N__21337\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21219\,
            in2 => \_gnd_net_\,
            in3 => \N__21255\,
            lcout => \current_shift_inst.PI_CTRL.N_155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21287\,
            in1 => \N__21478\,
            in2 => \N__21497\,
            in3 => \N__21578\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21527\,
            in1 => \N__21395\,
            in2 => \N__21515\,
            in3 => \N__21382\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPN72_22_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21493\,
            in2 => \_gnd_net_\,
            in3 => \N__21541\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21286\,
            in1 => \N__21577\,
            in2 => \N__21383\,
            in3 => \N__21394\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21511\,
            in1 => \N__21526\,
            in2 => \N__21727\,
            in3 => \N__21559\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21430\,
            in1 => \N__21004\,
            in2 => \N__20579\,
            in3 => \N__20576\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_9_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__24438\,
            in1 => \N__25996\,
            in2 => \N__24752\,
            in3 => \N__21869\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44911\,
            ce => \N__25649\,
            sr => \N__44179\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_16_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001110"
        )
    port map (
            in0 => \N__24737\,
            in1 => \N__23340\,
            in2 => \N__26034\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44911\,
            ce => \N__25649\,
            sr => \N__44179\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_10_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__24741\,
            in1 => \N__21856\,
            in2 => \N__21833\,
            in3 => \N__25997\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44911\,
            ce => \N__25649\,
            sr => \N__44179\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_11_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__26003\,
            in1 => \N__24743\,
            in2 => \N__21831\,
            in3 => \N__21782\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44911\,
            ce => \N__25649\,
            sr => \N__44179\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_12_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21830\,
            in1 => \N__24738\,
            in2 => \N__20660\,
            in3 => \N__25998\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44911\,
            ce => \N__25649\,
            sr => \N__44179\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_13_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__26004\,
            in1 => \N__24744\,
            in2 => \N__21832\,
            in3 => \N__20633\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44911\,
            ce => \N__25649\,
            sr => \N__44179\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_15_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24742\,
            in1 => \N__25999\,
            in2 => \N__24893\,
            in3 => \N__24408\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44911\,
            ce => \N__25649\,
            sr => \N__44179\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_7_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__25523\,
            in1 => \_gnd_net_\,
            in2 => \N__26033\,
            in3 => \N__25805\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44911\,
            ce => \N__25649\,
            sr => \N__44179\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001110"
        )
    port map (
            in0 => \N__21896\,
            in1 => \N__31638\,
            in2 => \N__31864\,
            in3 => \N__22070\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__21929\,
            in1 => \N__22040\,
            in2 => \N__31649\,
            in3 => \N__31847\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101100"
        )
    port map (
            in0 => \N__22100\,
            in1 => \N__31637\,
            in2 => \N__31863\,
            in3 => \N__23336\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20600\,
            in3 => \N__25463\,
            lcout => \elapsed_time_ns_1_RNI3VBED1_0_16\,
            ltout => \elapsed_time_ns_1_RNI3VBED1_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_9_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__24464\,
            in1 => \N__23412\,
            in2 => \N__20597\,
            in3 => \N__23376\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_i_a2_10_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__21930\,
            in1 => \_gnd_net_\,
            in2 => \N__20594\,
            in3 => \N__24887\,
            lcout => \phase_controller_inst1.stoper_hc.N_315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__26339\,
            in1 => \N__31817\,
            in2 => \N__20774\,
            in3 => \N__20628\,
            lcout => \elapsed_time_ns_1_RNIQ2MD11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__31818\,
            in1 => \N__26340\,
            in2 => \N__20798\,
            in3 => \N__20653\,
            lcout => \elapsed_time_ns_1_RNIP1MD11_0_12\,
            ltout => \elapsed_time_ns_1_RNIP1MD11_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_12_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__24739\,
            in1 => \N__26038\,
            in2 => \N__20663\,
            in3 => \N__21824\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44903\,
            ce => \N__31528\,
            sr => \N__44188\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__31819\,
            in1 => \N__26341\,
            in2 => \N__20825\,
            in3 => \N__21777\,
            lcout => \elapsed_time_ns_1_RNIO0MD11_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__26338\,
            in1 => \N__31816\,
            in2 => \N__20846\,
            in3 => \N__21849\,
            lcout => \elapsed_time_ns_1_RNINVLD11_0_10\,
            ltout => \elapsed_time_ns_1_RNINVLD11_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2_2_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20624\,
            in1 => \N__20652\,
            in2 => \N__20639\,
            in3 => \N__21776\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a0_6_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__21888\,
            in1 => \_gnd_net_\,
            in2 => \N__20636\,
            in3 => \N__24883\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a5_1_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_13_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21823\,
            in1 => \N__24740\,
            in2 => \N__20632\,
            in3 => \N__26039\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44903\,
            ce => \N__31528\,
            sr => \N__44188\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20606\,
            in2 => \_gnd_net_\,
            in3 => \N__25449\,
            lcout => \elapsed_time_ns_1_RNI51CED1_0_18\,
            ltout => \elapsed_time_ns_1_RNI51CED1_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011011100"
        )
    port map (
            in0 => \N__31777\,
            in1 => \N__31621\,
            in2 => \N__20609\,
            in3 => \N__22121\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__23786\,
            in1 => \N__22069\,
            in2 => \N__22004\,
            in3 => \N__21956\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__31775\,
            in1 => \N__21758\,
            in2 => \N__20900\,
            in3 => \N__26331\,
            lcout => \elapsed_time_ns_1_RNIR4ND11_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__26332\,
            in1 => \N__31778\,
            in2 => \N__20744\,
            in3 => \N__24882\,
            lcout => \elapsed_time_ns_1_RNIS4MD11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__25450\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20684\,
            lcout => \elapsed_time_ns_1_RNIL13KD1_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__21746\,
            in1 => \N__20876\,
            in2 => \N__26373\,
            in3 => \N__31776\,
            lcout => \elapsed_time_ns_1_RNIS5ND11_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31570\,
            in1 => \N__22120\,
            in2 => \N__22099\,
            in3 => \N__22035\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23275\,
            in1 => \N__20893\,
            in2 => \N__23465\,
            in3 => \N__23224\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__25537\,
            in1 => \N__22061\,
            in2 => \_gnd_net_\,
            in3 => \N__24805\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__22036\,
            in1 => \N__20711\,
            in2 => \N__20675\,
            in3 => \N__20740\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__23527\,
            in1 => \N__23554\,
            in2 => \_gnd_net_\,
            in3 => \N__23497\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20872\,
            in1 => \N__23590\,
            in2 => \N__20672\,
            in3 => \N__20669\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20794\,
            in1 => \N__20818\,
            in2 => \N__20773\,
            in3 => \N__20839\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24804\,
            in1 => \N__25536\,
            in2 => \N__20705\,
            in3 => \N__20739\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22242\,
            in2 => \N__23696\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_7_18_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__44886\,
            ce => \N__23653\,
            sr => \N__44219\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22218\,
            in2 => \N__23675\,
            in3 => \N__20702\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__44886\,
            ce => \N__23653\,
            sr => \N__44219\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22194\,
            in2 => \N__22247\,
            in3 => \N__20699\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__44886\,
            ce => \N__23653\,
            sr => \N__44219\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22563\,
            in2 => \N__22223\,
            in3 => \N__20696\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__44886\,
            ce => \N__23653\,
            sr => \N__44219\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22542\,
            in2 => \N__22199\,
            in3 => \N__20693\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__44886\,
            ce => \N__23653\,
            sr => \N__44219\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22524\,
            in2 => \N__22568\,
            in3 => \N__20690\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__44886\,
            ce => \N__23653\,
            sr => \N__44219\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22543\,
            in2 => \N__22508\,
            in3 => \N__20687\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__44886\,
            ce => \N__23653\,
            sr => \N__44219\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22525\,
            in2 => \N__22475\,
            in3 => \N__20828\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__44886\,
            ce => \N__23653\,
            sr => \N__44219\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22440\,
            in2 => \N__22504\,
            in3 => \N__20801\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__44878\,
            ce => \N__23652\,
            sr => \N__44225\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22416\,
            in2 => \N__22474\,
            in3 => \N__20777\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__44878\,
            ce => \N__23652\,
            sr => \N__44225\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22392\,
            in2 => \N__22445\,
            in3 => \N__20750\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__44878\,
            ce => \N__23652\,
            sr => \N__44225\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22755\,
            in2 => \N__22421\,
            in3 => \N__20747\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__44878\,
            ce => \N__23652\,
            sr => \N__44225\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22734\,
            in2 => \N__22397\,
            in3 => \N__20723\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__44878\,
            ce => \N__23652\,
            sr => \N__44225\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22716\,
            in2 => \N__22760\,
            in3 => \N__20720\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__44878\,
            ce => \N__23652\,
            sr => \N__44225\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22735\,
            in2 => \N__22700\,
            in3 => \N__20717\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__44878\,
            ce => \N__23652\,
            sr => \N__44225\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22717\,
            in2 => \N__22670\,
            in3 => \N__20714\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__44878\,
            ce => \N__23652\,
            sr => \N__44225\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22635\,
            in2 => \N__22699\,
            in3 => \N__20912\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__44872\,
            ce => \N__23651\,
            sr => \N__44230\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22611\,
            in2 => \N__22669\,
            in3 => \N__20909\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__44872\,
            ce => \N__23651\,
            sr => \N__44230\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22587\,
            in2 => \N__22640\,
            in3 => \N__20906\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__44872\,
            ce => \N__23651\,
            sr => \N__44230\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22953\,
            in2 => \N__22616\,
            in3 => \N__20903\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__44872\,
            ce => \N__23651\,
            sr => \N__44230\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22932\,
            in2 => \N__22592\,
            in3 => \N__20879\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__44872\,
            ce => \N__23651\,
            sr => \N__44230\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22914\,
            in2 => \N__22958\,
            in3 => \N__20858\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__44872\,
            ce => \N__23651\,
            sr => \N__44230\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22933\,
            in2 => \N__22898\,
            in3 => \N__20855\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__44872\,
            ce => \N__23651\,
            sr => \N__44230\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22915\,
            in2 => \N__22868\,
            in3 => \N__20852\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__44872\,
            ce => \N__23651\,
            sr => \N__44230\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22833\,
            in2 => \N__22897\,
            in3 => \N__20849\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__44865\,
            ce => \N__23650\,
            sr => \N__44233\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22809\,
            in2 => \N__22867\,
            in3 => \N__20990\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__44865\,
            ce => \N__23650\,
            sr => \N__44233\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22789\,
            in2 => \N__22838\,
            in3 => \N__20987\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__44865\,
            ce => \N__23650\,
            sr => \N__44233\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22771\,
            in2 => \N__22814\,
            in3 => \N__20984\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__44865\,
            ce => \N__23650\,
            sr => \N__44233\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20981\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44865\,
            ce => \N__23650\,
            sr => \N__44233\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20978\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23069\,
            in2 => \N__32414\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__44921\,
            ce => 'H',
            sr => \N__44152\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25028\,
            in2 => \N__32345\,
            in3 => \N__20933\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__44921\,
            ce => 'H',
            sr => \N__44152\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34490\,
            in2 => \N__23108\,
            in3 => \N__20915\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__44921\,
            ce => 'H',
            sr => \N__44152\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23090\,
            in2 => \N__32255\,
            in3 => \N__21242\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__44921\,
            ce => 'H',
            sr => \N__44152\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30302\,
            in2 => \N__23099\,
            in3 => \N__21203\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__44921\,
            ce => 'H',
            sr => \N__44152\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31268\,
            in2 => \N__23084\,
            in3 => \N__21167\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__44921\,
            ce => 'H',
            sr => \N__44152\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23882\,
            in2 => \N__34649\,
            in3 => \N__21131\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__44921\,
            ce => 'H',
            sr => \N__44152\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23075\,
            in2 => \N__30647\,
            in3 => \N__21098\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__44921\,
            ce => 'H',
            sr => \N__44152\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25274\,
            in2 => \N__30443\,
            in3 => \N__21056\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__44915\,
            ce => 'H',
            sr => \N__44159\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23873\,
            in2 => \N__31100\,
            in3 => \N__21023\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__44915\,
            ce => 'H',
            sr => \N__44159\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25265\,
            in2 => \N__35333\,
            in3 => \N__21011\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__44915\,
            ce => 'H',
            sr => \N__44159\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23063\,
            in2 => \N__34232\,
            in3 => \N__20993\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__44915\,
            ce => 'H',
            sr => \N__44159\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22994\,
            in2 => \N__30536\,
            in3 => \N__21398\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__44915\,
            ce => 'H',
            sr => \N__44159\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30907\,
            in2 => \N__23035\,
            in3 => \N__21386\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__44915\,
            ce => 'H',
            sr => \N__44159\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22998\,
            in2 => \N__34397\,
            in3 => \N__21368\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__44915\,
            ce => 'H',
            sr => \N__44159\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30383\,
            in2 => \N__23036\,
            in3 => \N__21347\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__44915\,
            ce => 'H',
            sr => \N__44159\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30809\,
            in2 => \N__23037\,
            in3 => \N__21326\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__44912\,
            ce => 'H',
            sr => \N__44164\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23005\,
            in2 => \N__31013\,
            in3 => \N__21311\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__44912\,
            ce => 'H',
            sr => \N__44164\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30707\,
            in2 => \N__23038\,
            in3 => \N__21290\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__44912\,
            ce => 'H',
            sr => \N__44164\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23009\,
            in2 => \N__34346\,
            in3 => \N__21278\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__44912\,
            ce => 'H',
            sr => \N__44164\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32618\,
            in2 => \N__23039\,
            in3 => \N__21569\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__44912\,
            ce => 'H',
            sr => \N__44164\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23013\,
            in2 => \N__32564\,
            in3 => \N__21548\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__44912\,
            ce => 'H',
            sr => \N__44164\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32510\,
            in2 => \N__23040\,
            in3 => \N__21530\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__44912\,
            ce => 'H',
            sr => \N__44164\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23017\,
            in2 => \N__35228\,
            in3 => \N__21518\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__44912\,
            ce => 'H',
            sr => \N__44164\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23041\,
            in2 => \N__35171\,
            in3 => \N__21500\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__44908\,
            ce => 'H',
            sr => \N__44174\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35111\,
            in2 => \N__23055\,
            in3 => \N__21485\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__44908\,
            ce => 'H',
            sr => \N__44174\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23045\,
            in2 => \N__35054\,
            in3 => \N__21464\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__44908\,
            ce => 'H',
            sr => \N__44174\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28664\,
            in2 => \N__23056\,
            in3 => \N__21440\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__44908\,
            ce => 'H',
            sr => \N__44174\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23049\,
            in2 => \N__34595\,
            in3 => \N__21419\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__44908\,
            ce => 'H',
            sr => \N__44174\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34532\,
            in2 => \N__23057\,
            in3 => \N__21707\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__44908\,
            ce => 'H',
            sr => \N__44174\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23053\,
            in2 => \N__35885\,
            in3 => \N__21683\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__44908\,
            ce => 'H',
            sr => \N__44174\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23054\,
            in1 => \N__35834\,
            in2 => \_gnd_net_\,
            in3 => \N__21680\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44908\,
            ce => 'H',
            sr => \N__44174\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_14_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24891\,
            in2 => \_gnd_net_\,
            in3 => \N__24404\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25256\,
            in2 => \_gnd_net_\,
            in3 => \N__25202\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_i_1_9_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__21895\,
            in1 => \N__24701\,
            in2 => \_gnd_net_\,
            in3 => \N__21816\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__31854\,
            in1 => \N__23416\,
            in2 => \N__31650\,
            in3 => \N__22151\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__24542\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25464\,
            lcout => \elapsed_time_ns_1_RNI62CED1_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_14_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__21934\,
            in1 => \N__21589\,
            in2 => \N__24727\,
            in3 => \N__26010\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44897\,
            ce => \N__31527\,
            sr => \N__44184\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_9_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__26011\,
            in1 => \N__21868\,
            in2 => \N__24439\,
            in3 => \N__24699\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44897\,
            ce => \N__31527\,
            sr => \N__44184\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_15_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__24881\,
            in1 => \N__26015\,
            in2 => \N__24726\,
            in3 => \N__24409\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44897\,
            ce => \N__31527\,
            sr => \N__44184\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_18_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001110"
        )
    port map (
            in0 => \N__23375\,
            in1 => \N__24691\,
            in2 => \N__26037\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44897\,
            ce => \N__31527\,
            sr => \N__44184\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_17_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__24688\,
            in1 => \N__26008\,
            in2 => \_gnd_net_\,
            in3 => \N__23411\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44897\,
            ce => \N__31527\,
            sr => \N__44184\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_16_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001110"
        )
    port map (
            in0 => \N__23341\,
            in1 => \N__24690\,
            in2 => \N__26036\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44897\,
            ce => \N__31527\,
            sr => \N__44184\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_10_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__24689\,
            in1 => \N__26009\,
            in2 => \N__21857\,
            in3 => \N__21826\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44897\,
            ce => \N__31527\,
            sr => \N__44184\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_11_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__21825\,
            in1 => \N__24692\,
            in2 => \N__26035\,
            in3 => \N__21781\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44897\,
            ce => \N__31527\,
            sr => \N__44184\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_i_o5_0_15_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21757\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21745\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_i_o5_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__44321\,
            in1 => \N__22340\,
            in2 => \N__22325\,
            in3 => \N__23739\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__44326\,
            in1 => \N__24522\,
            in2 => \N__21977\,
            in3 => \N__21986\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__21974\,
            in1 => \_gnd_net_\,
            in2 => \N__21965\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNI40CED1_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1_6_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21922\,
            in2 => \_gnd_net_\,
            in3 => \N__24868\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__24523\,
            in1 => \N__22276\,
            in2 => \N__44338\,
            in3 => \N__23771\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__23740\,
            in1 => \N__44322\,
            in2 => \N__21962\,
            in3 => \N__22175\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__26120\,
            in1 => \N__31808\,
            in2 => \N__21959\,
            in3 => \N__22361\,
            lcout => \elapsed_time_ns_1_RNIB4DJ11_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23712\,
            in2 => \_gnd_net_\,
            in3 => \N__26248\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25448\,
            in2 => \_gnd_net_\,
            in3 => \N__21950\,
            lcout => \elapsed_time_ns_1_RNI1TBED1_0_14\,
            ltout => \elapsed_time_ns_1_RNI1TBED1_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_9_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24864\,
            in2 => \N__21899\,
            in3 => \N__21887\,
            lcout => \phase_controller_inst1.stoper_hc.N_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44331\,
            in1 => \N__24526\,
            in2 => \_gnd_net_\,
            in3 => \N__22294\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24571\,
            in1 => \N__22150\,
            in2 => \N__22169\,
            in3 => \N__22160\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22154\,
            in3 => \N__23752\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_382_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__23299\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23197\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__25368\,
            in1 => \N__31809\,
            in2 => \N__26394\,
            in3 => \N__22373\,
            lcout => \elapsed_time_ns_1_RNIA3DJ11_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22137\,
            in1 => \N__22114\,
            in2 => \N__22098\,
            in3 => \N__24564\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22065\,
            in1 => \N__22034\,
            in2 => \N__22010\,
            in3 => \N__31566\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22317\,
            in1 => \N__44333\,
            in2 => \N__22007\,
            in3 => \N__22003\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__22339\,
            in1 => \_gnd_net_\,
            in2 => \N__21989\,
            in3 => \N__23766\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22372\,
            in2 => \_gnd_net_\,
            in3 => \N__22357\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__22298\,
            in1 => \N__24525\,
            in2 => \N__22280\,
            in3 => \N__23767\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111001111"
        )
    port map (
            in0 => \N__22346\,
            in1 => \N__22338\,
            in2 => \N__22324\,
            in3 => \N__22304\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24524\,
            in2 => \N__22283\,
            in3 => \N__22269\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29030\,
            in1 => \N__23691\,
            in2 => \_gnd_net_\,
            in3 => \N__22253\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__44873\,
            ce => \N__25595\,
            sr => \N__44220\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29003\,
            in1 => \N__23670\,
            in2 => \_gnd_net_\,
            in3 => \N__22250\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__44873\,
            ce => \N__25595\,
            sr => \N__44220\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29031\,
            in1 => \N__22243\,
            in2 => \_gnd_net_\,
            in3 => \N__22226\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__44873\,
            ce => \N__25595\,
            sr => \N__44220\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29004\,
            in1 => \N__22219\,
            in2 => \_gnd_net_\,
            in3 => \N__22202\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__44873\,
            ce => \N__25595\,
            sr => \N__44220\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29032\,
            in1 => \N__22195\,
            in2 => \_gnd_net_\,
            in3 => \N__22178\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__44873\,
            ce => \N__25595\,
            sr => \N__44220\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29005\,
            in1 => \N__22564\,
            in2 => \_gnd_net_\,
            in3 => \N__22547\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__44873\,
            ce => \N__25595\,
            sr => \N__44220\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29033\,
            in1 => \N__22544\,
            in2 => \_gnd_net_\,
            in3 => \N__22529\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__44873\,
            ce => \N__25595\,
            sr => \N__44220\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29006\,
            in1 => \N__22526\,
            in2 => \_gnd_net_\,
            in3 => \N__22511\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__44873\,
            ce => \N__25595\,
            sr => \N__44220\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28977\,
            in1 => \N__22497\,
            in2 => \_gnd_net_\,
            in3 => \N__22478\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__44866\,
            ce => \N__25596\,
            sr => \N__44226\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29002\,
            in1 => \N__22467\,
            in2 => \_gnd_net_\,
            in3 => \N__22448\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__44866\,
            ce => \N__25596\,
            sr => \N__44226\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28974\,
            in1 => \N__22441\,
            in2 => \_gnd_net_\,
            in3 => \N__22424\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__44866\,
            ce => \N__25596\,
            sr => \N__44226\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28999\,
            in1 => \N__22417\,
            in2 => \_gnd_net_\,
            in3 => \N__22400\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__44866\,
            ce => \N__25596\,
            sr => \N__44226\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28975\,
            in1 => \N__22393\,
            in2 => \_gnd_net_\,
            in3 => \N__22376\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__44866\,
            ce => \N__25596\,
            sr => \N__44226\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29000\,
            in1 => \N__22756\,
            in2 => \_gnd_net_\,
            in3 => \N__22739\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__44866\,
            ce => \N__25596\,
            sr => \N__44226\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28976\,
            in1 => \N__22736\,
            in2 => \_gnd_net_\,
            in3 => \N__22721\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__44866\,
            ce => \N__25596\,
            sr => \N__44226\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29001\,
            in1 => \N__22718\,
            in2 => \_gnd_net_\,
            in3 => \N__22703\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__44866\,
            ce => \N__25596\,
            sr => \N__44226\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29007\,
            in1 => \N__22692\,
            in2 => \_gnd_net_\,
            in3 => \N__22673\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__44859\,
            ce => \N__25607\,
            sr => \N__44231\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29013\,
            in1 => \N__22662\,
            in2 => \_gnd_net_\,
            in3 => \N__22643\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__44859\,
            ce => \N__25607\,
            sr => \N__44231\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29008\,
            in1 => \N__22636\,
            in2 => \_gnd_net_\,
            in3 => \N__22619\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__44859\,
            ce => \N__25607\,
            sr => \N__44231\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29014\,
            in1 => \N__22612\,
            in2 => \_gnd_net_\,
            in3 => \N__22595\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__44859\,
            ce => \N__25607\,
            sr => \N__44231\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29009\,
            in1 => \N__22588\,
            in2 => \_gnd_net_\,
            in3 => \N__22571\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__44859\,
            ce => \N__25607\,
            sr => \N__44231\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29015\,
            in1 => \N__22954\,
            in2 => \_gnd_net_\,
            in3 => \N__22937\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__44859\,
            ce => \N__25607\,
            sr => \N__44231\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29010\,
            in1 => \N__22934\,
            in2 => \_gnd_net_\,
            in3 => \N__22919\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__44859\,
            ce => \N__25607\,
            sr => \N__44231\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29016\,
            in1 => \N__22916\,
            in2 => \_gnd_net_\,
            in3 => \N__22901\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__44859\,
            ce => \N__25607\,
            sr => \N__44231\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29017\,
            in1 => \N__22890\,
            in2 => \_gnd_net_\,
            in3 => \N__22871\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__44856\,
            ce => \N__25606\,
            sr => \N__44234\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29011\,
            in1 => \N__22860\,
            in2 => \_gnd_net_\,
            in3 => \N__22841\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__44856\,
            ce => \N__25606\,
            sr => \N__44234\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29018\,
            in1 => \N__22834\,
            in2 => \_gnd_net_\,
            in3 => \N__22817\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__44856\,
            ce => \N__25606\,
            sr => \N__44234\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29012\,
            in1 => \N__22810\,
            in2 => \_gnd_net_\,
            in3 => \N__22793\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__44856\,
            ce => \N__25606\,
            sr => \N__44234\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29019\,
            in1 => \N__22790\,
            in2 => \_gnd_net_\,
            in3 => \N__22778\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__44856\,
            ce => \N__25606\,
            sr => \N__44234\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__22772\,
            in1 => \N__29020\,
            in2 => \_gnd_net_\,
            in3 => \N__22775\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44856\,
            ce => \N__25606\,
            sr => \N__44234\
        );

    \phase_controller_inst2.S2_LC_8_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26603\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44833\,
            ce => 'H',
            sr => \N__44239\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28427\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44916\,
            ce => 'H',
            sr => \N__44146\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28277\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44916\,
            ce => 'H',
            sr => \N__44146\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28400\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44916\,
            ce => 'H',
            sr => \N__44146\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26909\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44916\,
            ce => 'H',
            sr => \N__44146\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28298\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44916\,
            ce => 'H',
            sr => \N__44146\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28256\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44913\,
            ce => 'H',
            sr => \N__44153\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30250\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44913\,
            ce => 'H',
            sr => \N__44153\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34942\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44913\,
            ce => 'H',
            sr => \N__44153\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23144\,
            in2 => \N__25157\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23828\,
            in2 => \_gnd_net_\,
            in3 => \N__23138\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \N__44904\,
            ce => 'H',
            sr => \N__25130\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23807\,
            in2 => \N__25016\,
            in3 => \N__23135\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \N__44904\,
            ce => 'H',
            sr => \N__25130\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24134\,
            in2 => \_gnd_net_\,
            in3 => \N__23132\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \N__44904\,
            ce => 'H',
            sr => \N__25130\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24110\,
            in2 => \_gnd_net_\,
            in3 => \N__23129\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \N__44904\,
            ce => 'H',
            sr => \N__25130\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24086\,
            in2 => \_gnd_net_\,
            in3 => \N__23126\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \N__44904\,
            ce => 'H',
            sr => \N__25130\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24050\,
            in2 => \_gnd_net_\,
            in3 => \N__23123\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \N__44904\,
            ce => 'H',
            sr => \N__25130\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24029\,
            in2 => \_gnd_net_\,
            in3 => \N__23120\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \N__44904\,
            ce => 'H',
            sr => \N__25130\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23993\,
            in2 => \_gnd_net_\,
            in3 => \N__23117\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \N__44898\,
            ce => 'H',
            sr => \N__25126\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23960\,
            in2 => \_gnd_net_\,
            in3 => \N__23171\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \N__44898\,
            ce => 'H',
            sr => \N__25126\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23939\,
            in2 => \_gnd_net_\,
            in3 => \N__23168\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \N__44898\,
            ce => 'H',
            sr => \N__25126\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24374\,
            in2 => \_gnd_net_\,
            in3 => \N__23165\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \N__44898\,
            ce => 'H',
            sr => \N__25126\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24326\,
            in2 => \_gnd_net_\,
            in3 => \N__23162\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \N__44898\,
            ce => 'H',
            sr => \N__25126\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24305\,
            in2 => \_gnd_net_\,
            in3 => \N__23159\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \N__44898\,
            ce => 'H',
            sr => \N__25126\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24263\,
            in2 => \_gnd_net_\,
            in3 => \N__23156\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \N__44898\,
            ce => 'H',
            sr => \N__25126\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24230\,
            in2 => \_gnd_net_\,
            in3 => \N__23153\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \N__44898\,
            ce => 'H',
            sr => \N__25126\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24191\,
            in2 => \_gnd_net_\,
            in3 => \N__23150\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \N__44892\,
            ce => 'H',
            sr => \N__25118\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24155\,
            in2 => \_gnd_net_\,
            in3 => \N__23147\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \N__44892\,
            ce => 'H',
            sr => \N__25118\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24605\,
            in2 => \_gnd_net_\,
            in3 => \N__23423\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44892\,
            ce => 'H',
            sr => \N__25118\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3_2_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23401\,
            in1 => \N__25361\,
            in2 => \N__26121\,
            in3 => \N__23377\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_2_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24474\,
            in1 => \N__23345\,
            in2 => \N__23315\,
            in3 => \N__23312\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__31802\,
            in1 => \N__23252\,
            in2 => \N__26381\,
            in3 => \N__23306\,
            lcout => \elapsed_time_ns_1_RNIP2ND11_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__23258\,
            in1 => \N__26348\,
            in2 => \N__23285\,
            in3 => \N__31801\,
            lcout => \elapsed_time_ns_1_RNI1BND11_0_29\,
            ltout => \elapsed_time_ns_1_RNI1BND11_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_i_o5_7_15_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23438\,
            in1 => \N__23251\,
            in2 => \N__23243\,
            in3 => \N__23209\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_7_i_o5_7Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_i_o5_15_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23240\,
            in1 => \N__23179\,
            in2 => \N__23234\,
            in3 => \N__23561\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__31803\,
            in1 => \N__23210\,
            in2 => \N__26382\,
            in3 => \N__23231\,
            lcout => \elapsed_time_ns_1_RNIO1ND11_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__23201\,
            in1 => \N__23180\,
            in2 => \N__26398\,
            in3 => \N__31804\,
            lcout => \elapsed_time_ns_1_RNIQ3ND11_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_4_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__25939\,
            in1 => \N__25799\,
            in2 => \N__25372\,
            in3 => \N__25728\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44879\,
            ce => \N__31529\,
            sr => \N__44189\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__26333\,
            in1 => \N__31771\,
            in2 => \N__23573\,
            in3 => \N__23594\,
            lcout => \elapsed_time_ns_1_RNIT6ND11_0_25\,
            ltout => \elapsed_time_ns_1_RNIT6ND11_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_i_o5_6_15_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23476\,
            in1 => \N__23536\,
            in2 => \N__23564\,
            in3 => \N__23509\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_i_o5_6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__23537\,
            in1 => \N__23555\,
            in2 => \N__26374\,
            in3 => \N__31774\,
            lcout => \elapsed_time_ns_1_RNIV8ND11_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__31772\,
            in1 => \N__23528\,
            in2 => \N__26396\,
            in3 => \N__23510\,
            lcout => \elapsed_time_ns_1_RNIU7ND11_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__26334\,
            in1 => \N__23501\,
            in2 => \N__23480\,
            in3 => \N__31773\,
            lcout => \elapsed_time_ns_1_RNI0AND11_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_5_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__25940\,
            in1 => \N__25800\,
            in2 => \N__26125\,
            in3 => \N__25729\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44879\,
            ce => \N__31529\,
            sr => \N__44189\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__31799\,
            in1 => \N__23464\,
            in2 => \N__26395\,
            in3 => \N__23437\,
            lcout => \elapsed_time_ns_1_RNIP3OD11_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23785\,
            in1 => \N__25486\,
            in2 => \N__23723\,
            in3 => \N__26244\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__44332\,
            in1 => \N__23753\,
            in2 => \_gnd_net_\,
            in3 => \N__23741\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__26204\,
            in1 => \N__31800\,
            in2 => \N__23726\,
            in3 => \N__23722\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23699\,
            in3 => \N__31608\,
            lcout => \elapsed_time_ns_1_RNIQURR91_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23695\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44867\,
            ce => \N__23654\,
            sr => \N__44210\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23674\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44867\,
            ce => \N__23654\,
            sr => \N__44210\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29065\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29104\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_432_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_1_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27895\,
            in2 => \_gnd_net_\,
            in3 => \N__24927\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23612\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S1_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27907\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44836\,
            ce => 'H',
            sr => \N__44238\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23897\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34453\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44909\,
            ce => 'H',
            sr => \N__44135\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31226\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44905\,
            ce => 'H',
            sr => \N__44143\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23864\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44899\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23855\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44899\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25817\,
            in2 => \N__23837\,
            in3 => \N__25146\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25388\,
            in2 => \N__23816\,
            in3 => \N__23827\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23806\,
            in1 => \N__25661\,
            in2 => \N__23795\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24133\,
            in1 => \N__25340\,
            in2 => \N__24122\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26090\,
            in2 => \N__24098\,
            in3 => \N__24109\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24085\,
            in1 => \N__25415\,
            in2 => \N__24074\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24062\,
            in2 => \N__24038\,
            in3 => \N__24049\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26051\,
            in2 => \N__24017\,
            in3 => \N__24028\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24005\,
            in2 => \N__23981\,
            in3 => \N__23992\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23972\,
            in2 => \N__23948\,
            in3 => \N__23959\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23938\,
            in1 => \N__23927\,
            in2 => \N__23915\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24373\,
            in1 => \N__24362\,
            in2 => \N__24350\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24341\,
            in2 => \N__24314\,
            in3 => \N__24325\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24304\,
            in1 => \N__24281\,
            in2 => \N__24293\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24275\,
            in2 => \N__24251\,
            in3 => \N__24262\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24242\,
            in2 => \N__24218\,
            in3 => \N__24229\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24206\,
            in2 => \N__24179\,
            in3 => \N__24190\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24170\,
            in2 => \N__24143\,
            in3 => \N__24154\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24620\,
            in2 => \N__24593\,
            in3 => \N__24604\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24584\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__31859\,
            in1 => \N__24482\,
            in2 => \N__31658\,
            in3 => \N__24572\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__24530\,
            in1 => \N__26390\,
            in2 => \N__26022\,
            in3 => \N__31858\,
            lcout => \elapsed_time_ns_1_RNIQ4OD11_0_31\,
            ltout => \elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_19_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001110"
        )
    port map (
            in0 => \N__24674\,
            in1 => \N__24481\,
            in2 => \N__24443\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44874\,
            ce => \N__31526\,
            sr => \N__44175\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_3_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__25785\,
            in1 => \N__26209\,
            in2 => \N__25733\,
            in3 => \N__25673\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44874\,
            ce => \N__31526\,
            sr => \N__44175\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_0_6_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__24440\,
            in1 => \N__24413\,
            in2 => \N__24700\,
            in3 => \N__24383\,
            lcout => \phase_controller_inst1.stoper_hc.N_325\,
            ltout => \phase_controller_inst1.stoper_hc.N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_6_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__25981\,
            in1 => \N__31683\,
            in2 => \N__24908\,
            in3 => \N__25730\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44874\,
            ce => \N__31526\,
            sr => \N__44175\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0_2_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__25515\,
            in1 => \N__31679\,
            in2 => \N__26077\,
            in3 => \N__24905\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_6_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24892\,
            in2 => \N__24821\,
            in3 => \N__24668\,
            lcout => \phase_controller_inst1.stoper_hc.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_i_0_2_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__24771\,
            in1 => \N__26200\,
            in2 => \N__24791\,
            in3 => \N__26225\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_i_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_0_a5_1_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__24786\,
            in1 => \N__26171\,
            in2 => \N__24772\,
            in3 => \N__24669\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.N_307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_0_1_1_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25714\,
            in2 => \N__24818\,
            in3 => \N__25845\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_f0_0_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__31835\,
            in1 => \N__26399\,
            in2 => \N__24815\,
            in3 => \N__26072\,
            lcout => \elapsed_time_ns_1_RNIE7DJ11_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31547\,
            in2 => \_gnd_net_\,
            in3 => \N__25472\,
            lcout => \elapsed_time_ns_1_RNIIU2KD1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_0_0_3_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__24787\,
            in1 => \N__25911\,
            in2 => \N__24773\,
            in3 => \N__24670\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_7_f0_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNI41671_0_1_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__24970\,
            in1 => \N__44327\,
            in2 => \N__25248\,
            in3 => \N__24996\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUB_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25234\,
            in2 => \_gnd_net_\,
            in3 => \N__25194\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000100010"
        )
    port map (
            in0 => \N__25239\,
            in1 => \N__25199\,
            in2 => \N__24977\,
            in3 => \N__24997\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44861\,
            ce => 'H',
            sr => \N__44185\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNI41671_1_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110110"
        )
    port map (
            in0 => \N__24994\,
            in1 => \N__24969\,
            in2 => \N__44339\,
            in3 => \N__25235\,
            lcout => \phase_controller_inst1.stoper_hc.un1_stoper_state12_1_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24971\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24995\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.N_45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__36623\,
            in1 => \N__25240\,
            in2 => \N__25001\,
            in3 => \N__25195\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44861\,
            ce => 'H',
            sr => \N__44185\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__24998\,
            in1 => \N__25244\,
            in2 => \N__24976\,
            in3 => \N__25200\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44857\,
            ce => 'H',
            sr => \N__44199\
        );

    \phase_controller_inst1.start_timer_hc_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__26665\,
            in1 => \N__26135\,
            in2 => \N__24975\,
            in3 => \N__36572\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44852\,
            ce => 'H',
            sr => \N__44208\
        );

    \phase_controller_inst2.state_2_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__24937\,
            in1 => \N__28011\,
            in2 => \N__27905\,
            in3 => \N__26447\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44848\,
            ce => 'H',
            sr => \N__44214\
        );

    \phase_controller_inst2.state_3_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__27891\,
            in1 => \N__28037\,
            in2 => \N__24938\,
            in3 => \N__25051\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44845\,
            ce => 'H',
            sr => \N__44221\
        );

    \phase_controller_inst2.T12_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__26590\,
            in1 => \N__28015\,
            in2 => \_gnd_net_\,
            in3 => \N__25063\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44845\,
            ce => 'H',
            sr => \N__44221\
        );

    \phase_controller_inst1.state_3_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__28838\,
            in1 => \N__25052\,
            in2 => \N__28895\,
            in3 => \N__26162\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44845\,
            ce => 'H',
            sr => \N__44221\
        );

    \phase_controller_inst2.state_ns_i_a3_1_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26701\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26650\,
            lcout => state_ns_i_a3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29135\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25042\,
            ce => 'H',
            sr => \N__44122\
        );

    \delay_measurement_inst.stop_timer_hc_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29136\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25043\,
            ce => 'H',
            sr => \N__44124\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30432\,
            in1 => \N__34644\,
            in2 => \N__31096\,
            in3 => \N__30643\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__30301\,
            in1 => \N__32247\,
            in2 => \N__25031\,
            in3 => \N__31263\,
            lcout => \current_shift_inst.PI_CTRL.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34528\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26797\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44900\,
            ce => 'H',
            sr => \N__44136\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28232\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44900\,
            ce => 'H',
            sr => \N__44136\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30334\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44900\,
            ce => 'H',
            sr => \N__44136\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34986\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44900\,
            ce => 'H',
            sr => \N__44136\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__25255\,
            in1 => \N__25201\,
            in2 => \_gnd_net_\,
            in3 => \N__25150\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44894\,
            ce => 'H',
            sr => \N__25125\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26483\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26824\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26423\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26525\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28709\,
            in2 => \N__25562\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27124\,
            in2 => \_gnd_net_\,
            in3 => \N__25079\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \N__44888\,
            ce => 'H',
            sr => \N__31409\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26924\,
            in2 => \N__27101\,
            in3 => \N__25301\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \N__44888\,
            ce => 'H',
            sr => \N__31409\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27049\,
            in2 => \_gnd_net_\,
            in3 => \N__25298\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \N__44888\,
            ce => 'H',
            sr => \N__31409\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27025\,
            in2 => \_gnd_net_\,
            in3 => \N__25295\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \N__44888\,
            ce => 'H',
            sr => \N__31409\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27445\,
            in2 => \_gnd_net_\,
            in3 => \N__25292\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \N__44888\,
            ce => 'H',
            sr => \N__31409\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27403\,
            in2 => \_gnd_net_\,
            in3 => \N__25289\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \N__44888\,
            ce => 'H',
            sr => \N__31409\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27376\,
            in2 => \_gnd_net_\,
            in3 => \N__25286\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \N__44888\,
            ce => 'H',
            sr => \N__31409\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27325\,
            in2 => \_gnd_net_\,
            in3 => \N__25283\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \N__44882\,
            ce => 'H',
            sr => \N__31408\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27289\,
            in2 => \_gnd_net_\,
            in3 => \N__25280\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \N__44882\,
            ce => 'H',
            sr => \N__31408\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27262\,
            in2 => \_gnd_net_\,
            in3 => \N__25277\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \N__44882\,
            ce => 'H',
            sr => \N__31408\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27211\,
            in2 => \_gnd_net_\,
            in3 => \N__25325\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \N__44882\,
            ce => 'H',
            sr => \N__31408\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27187\,
            in2 => \_gnd_net_\,
            in3 => \N__25322\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \N__44882\,
            ce => 'H',
            sr => \N__31408\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27679\,
            in2 => \_gnd_net_\,
            in3 => \N__25319\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \N__44882\,
            ce => 'H',
            sr => \N__31408\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27628\,
            in2 => \_gnd_net_\,
            in3 => \N__25316\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \N__44882\,
            ce => 'H',
            sr => \N__31408\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27601\,
            in2 => \_gnd_net_\,
            in3 => \N__25313\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \N__44882\,
            ce => 'H',
            sr => \N__31408\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27562\,
            in2 => \_gnd_net_\,
            in3 => \N__25310\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \N__44875\,
            ce => 'H',
            sr => \N__31400\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27526\,
            in2 => \_gnd_net_\,
            in3 => \N__25307\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \N__44875\,
            ce => 'H',
            sr => \N__31400\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27478\,
            in2 => \_gnd_net_\,
            in3 => \N__25304\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44875\,
            ce => 'H',
            sr => \N__31400\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_8_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25788\,
            in1 => \N__25931\,
            in2 => \_gnd_net_\,
            in3 => \N__26076\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44868\,
            ce => \N__31522\,
            sr => \N__44168\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__31855\,
            in1 => \N__26389\,
            in2 => \N__25547\,
            in3 => \N__25519\,
            lcout => \elapsed_time_ns_1_RNID6DJ11_0_7\,
            ltout => \elapsed_time_ns_1_RNID6DJ11_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_7_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__25787\,
            in1 => \_gnd_net_\,
            in2 => \N__25499\,
            in3 => \N__25932\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44868\,
            ce => \N__31522\,
            sr => \N__44168\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001110"
        )
    port map (
            in0 => \N__31856\,
            in1 => \N__31645\,
            in2 => \N__25496\,
            in3 => \N__25846\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25475\,
            in3 => \N__25468\,
            lcout => \elapsed_time_ns_1_RNIDP2KD1_0_1\,
            ltout => \elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_1_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__25929\,
            in1 => \N__25789\,
            in2 => \N__25418\,
            in3 => \N__25829\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44868\,
            ce => \N__31522\,
            sr => \N__44168\
        );

    \phase_controller_inst2.stoper_hc.target_time_esr_2_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__25786\,
            in1 => \N__25930\,
            in2 => \N__25732\,
            in3 => \N__25402\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44868\,
            ce => \N__31522\,
            sr => \N__44168\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_6_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__25720\,
            in1 => \N__25935\,
            in2 => \N__31687\,
            in3 => \N__25797\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44862\,
            ce => \N__25642\,
            sr => \N__44176\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_2_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__25937\,
            in1 => \N__25790\,
            in2 => \N__25403\,
            in3 => \N__25721\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44862\,
            ce => \N__25642\,
            sr => \N__44176\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_4_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__25719\,
            in1 => \N__25934\,
            in2 => \N__25376\,
            in3 => \N__25796\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44862\,
            ce => \N__25642\,
            sr => \N__44176\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_5_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__25938\,
            in1 => \N__25715\,
            in2 => \N__26129\,
            in3 => \N__25791\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44862\,
            ce => \N__25642\,
            sr => \N__44176\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_8_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25933\,
            in2 => \N__26078\,
            in3 => \N__25798\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44862\,
            ce => \N__25642\,
            sr => \N__44176\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_1_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__25936\,
            in1 => \N__25850\,
            in2 => \N__25804\,
            in3 => \N__25828\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44862\,
            ce => \N__25642\,
            sr => \N__44176\
        );

    \phase_controller_inst1.stoper_hc.target_time_esr_3_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__26210\,
            in1 => \N__25792\,
            in2 => \N__25731\,
            in3 => \N__25672\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44862\,
            ce => \N__25642\,
            sr => \N__44176\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40218\,
            in1 => \N__38435\,
            in2 => \_gnd_net_\,
            in3 => \N__38402\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__29066\,
            in1 => \N__29143\,
            in2 => \_gnd_net_\,
            in3 => \N__29097\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_433_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28559\,
            in2 => \_gnd_net_\,
            in3 => \N__28578\,
            lcout => \phase_controller_inst1.stoper_tr.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31458\,
            in2 => \_gnd_net_\,
            in3 => \N__28797\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26411\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__26397\,
            in1 => \N__31857\,
            in2 => \N__26255\,
            in3 => \N__26224\,
            lcout => \elapsed_time_ns_1_RNI81DJ11_0_2\,
            ltout => \elapsed_time_ns_1_RNI81DJ11_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_f0_0_o2_1_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26213\,
            in3 => \N__26205\,
            lcout => \phase_controller_inst1.stoper_hc.N_283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26501\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29413\,
            in2 => \_gnd_net_\,
            in3 => \N__28761\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__28579\,
            in1 => \N__26666\,
            in2 => \N__26165\,
            in3 => \N__26158\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44853\,
            ce => 'H',
            sr => \N__44186\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28732\,
            in2 => \_gnd_net_\,
            in3 => \N__26143\,
            lcout => \phase_controller_inst1.N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_0_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__29414\,
            in1 => \N__28762\,
            in2 => \N__26147\,
            in3 => \N__28733\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44853\,
            ce => 'H',
            sr => \N__44186\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28852\,
            in2 => \_gnd_net_\,
            in3 => \N__28890\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28009\,
            in2 => \_gnd_net_\,
            in3 => \N__26444\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.start_timer_hc_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__32007\,
            in1 => \N__26459\,
            in2 => \N__26450\,
            in3 => \N__26663\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44849\,
            ce => 'H',
            sr => \N__44200\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110001000"
        )
    port map (
            in0 => \N__26445\,
            in1 => \N__31985\,
            in2 => \N__28814\,
            in3 => \N__31472\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44849\,
            ce => 'H',
            sr => \N__44200\
        );

    \phase_controller_inst2.state_1_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__26623\,
            in1 => \N__28010\,
            in2 => \N__26592\,
            in3 => \N__26446\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44849\,
            ce => 'H',
            sr => \N__44200\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26580\,
            in2 => \_gnd_net_\,
            in3 => \N__26622\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.start_timer_tr_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__26664\,
            in1 => \N__43759\,
            in2 => \N__26429\,
            in3 => \N__28036\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44849\,
            ce => 'H',
            sr => \N__44200\
        );

    \current_shift_inst.control_input_0_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27728\,
            in2 => \N__39866\,
            in3 => \N__39864\,
            lcout => \current_shift_inst.control_inputZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \current_shift_inst.control_input_1_cry_0\,
            clk => \N__44846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27719\,
            in2 => \_gnd_net_\,
            in3 => \N__26426\,
            lcout => \current_shift_inst.control_inputZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_0\,
            carryout => \current_shift_inst.control_input_1_cry_1\,
            clk => \N__44846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_2_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27710\,
            in2 => \_gnd_net_\,
            in3 => \N__26414\,
            lcout => \current_shift_inst.control_inputZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_1\,
            carryout => \current_shift_inst.control_input_1_cry_2\,
            clk => \N__44846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_3_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27821\,
            in2 => \_gnd_net_\,
            in3 => \N__26402\,
            lcout => \current_shift_inst.control_inputZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_2\,
            carryout => \current_shift_inst.control_input_1_cry_3\,
            clk => \N__44846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_4_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27812\,
            in2 => \_gnd_net_\,
            in3 => \N__26510\,
            lcout => \current_shift_inst.control_inputZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_3\,
            carryout => \current_shift_inst.control_input_1_cry_4\,
            clk => \N__44846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_5_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27803\,
            in2 => \_gnd_net_\,
            in3 => \N__26507\,
            lcout => \current_shift_inst.control_inputZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_4\,
            carryout => \current_shift_inst.control_input_1_cry_5\,
            clk => \N__44846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_6_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27794\,
            in2 => \_gnd_net_\,
            in3 => \N__26504\,
            lcout => \current_shift_inst.control_inputZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_5\,
            carryout => \current_shift_inst.control_input_1_cry_6\,
            clk => \N__44846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_7_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27773\,
            in2 => \_gnd_net_\,
            in3 => \N__26492\,
            lcout => \current_shift_inst.control_inputZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_6\,
            carryout => \current_shift_inst.control_input_1_cry_7\,
            clk => \N__44846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_8_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27764\,
            in2 => \_gnd_net_\,
            in3 => \N__26489\,
            lcout => \current_shift_inst.control_inputZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \current_shift_inst.control_input_1_cry_8\,
            clk => \N__44843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_9_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27755\,
            in2 => \_gnd_net_\,
            in3 => \N__26486\,
            lcout => \current_shift_inst.control_inputZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_8\,
            carryout => \current_shift_inst.control_input_1_cry_9\,
            clk => \N__44843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_10_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26465\,
            in2 => \_gnd_net_\,
            in3 => \N__26471\,
            lcout => \current_shift_inst.control_inputZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_9\,
            carryout => \current_shift_inst.control_input_1_cry_10\,
            clk => \N__44843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_11_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001110111100010"
        )
    port map (
            in0 => \N__40125\,
            in1 => \N__28046\,
            in2 => \N__27743\,
            in3 => \N__26468\,
            lcout => \current_shift_inst.control_inputZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_c_RNIG7KU_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28045\,
            in2 => \_gnd_net_\,
            in3 => \N__27739\,
            lcout => \current_shift_inst.control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26729\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_4_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26700\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26651\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44841\,
            ce => 'H',
            sr => \N__44222\
        );

    \phase_controller_inst2.state_0_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__26627\,
            in1 => \N__40814\,
            in2 => \N__27938\,
            in3 => \N__26591\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44841\,
            ce => 'H',
            sr => \N__44222\
        );

    \phase_controller_inst2.T23_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__26536\,
            in1 => \N__26602\,
            in2 => \_gnd_net_\,
            in3 => \N__27936\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44839\,
            ce => 'H',
            sr => \N__44227\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31253\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30808\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31002\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30529\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34875\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35038\,
            in1 => \N__35099\,
            in2 => \N__34588\,
            in3 => \N__28661\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26741\,
            in1 => \N__30263\,
            in2 => \N__26744\,
            in3 => \N__28178\,
            lcout => \current_shift_inst.PI_CTRL.N_74_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32508\,
            in1 => \N__35166\,
            in2 => \N__32557\,
            in3 => \N__34342\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31341\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32246\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34882\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__30840\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34881\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30703\,
            in1 => \N__32612\,
            in2 => \N__31009\,
            in3 => \N__30382\,
            lcout => \current_shift_inst.PI_CTRL.N_74_16\,
            ltout => \current_shift_inst.PI_CTRL.N_74_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28147\,
            in1 => \N__28165\,
            in2 => \N__26732\,
            in3 => \N__34228\,
            lcout => \current_shift_inst.PI_CTRL.N_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__32338\,
            in1 => \N__34890\,
            in2 => \N__28352\,
            in3 => \N__26902\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34486\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34437\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32337\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26901\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34223\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26777\,
            in2 => \_gnd_net_\,
            in3 => \N__26801\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26933\,
            in2 => \_gnd_net_\,
            in3 => \N__26771\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__44893\,
            ce => 'H',
            sr => \N__44130\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26768\,
            in2 => \_gnd_net_\,
            in3 => \N__26762\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__44893\,
            ce => 'H',
            sr => \N__44130\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26759\,
            in2 => \_gnd_net_\,
            in3 => \N__26747\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__44893\,
            ce => 'H',
            sr => \N__44130\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26918\,
            in2 => \_gnd_net_\,
            in3 => \N__26912\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__44893\,
            ce => 'H',
            sr => \N__44130\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38327\,
            in2 => \_gnd_net_\,
            in3 => \N__26888\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__44893\,
            ce => 'H',
            sr => \N__44130\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26975\,
            in2 => \_gnd_net_\,
            in3 => \N__26885\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__44893\,
            ce => 'H',
            sr => \N__44130\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26882\,
            in2 => \_gnd_net_\,
            in3 => \N__26870\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__44893\,
            ce => 'H',
            sr => \N__44130\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26951\,
            in2 => \_gnd_net_\,
            in3 => \N__26867\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__44887\,
            ce => 'H',
            sr => \N__44137\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26864\,
            in2 => \_gnd_net_\,
            in3 => \N__26849\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__44887\,
            ce => 'H',
            sr => \N__44137\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26846\,
            in2 => \_gnd_net_\,
            in3 => \N__26840\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__44887\,
            ce => 'H',
            sr => \N__44137\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26837\,
            in2 => \_gnd_net_\,
            in3 => \N__26831\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__44887\,
            ce => 'H',
            sr => \N__44137\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26828\,
            in2 => \_gnd_net_\,
            in3 => \N__26804\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44887\,
            ce => 'H',
            sr => \N__44137\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__41880\,
            in1 => \N__43190\,
            in2 => \_gnd_net_\,
            in3 => \N__43148\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44880\,
            ce => 'H',
            sr => \N__39651\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26990\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26966\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30330\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31212\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26945\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHE_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31470\,
            in2 => \_gnd_net_\,
            in3 => \N__28809\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__31303\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34864\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34867\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31141\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__30594\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34865\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34866\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33268\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33526\,
            in2 => \_gnd_net_\,
            in3 => \N__34868\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28701\,
            in1 => \N__27149\,
            in2 => \N__27143\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27110\,
            in2 => \N__27134\,
            in3 => \N__27125\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27100\,
            in1 => \N__27068\,
            in2 => \N__27083\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27062\,
            in2 => \N__27035\,
            in3 => \N__27050\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27026\,
            in1 => \N__27011\,
            in2 => \N__26999\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27449\,
            in1 => \N__27431\,
            in2 => \N__27419\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27410\,
            in2 => \N__27389\,
            in3 => \N__27404\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27377\,
            in1 => \N__27362\,
            in2 => \N__27356\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27344\,
            in2 => \N__27311\,
            in3 => \N__27332\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27302\,
            in2 => \N__27275\,
            in3 => \N__27290\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27266\,
            in1 => \N__27248\,
            in2 => \N__27236\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27227\,
            in2 => \N__27197\,
            in3 => \N__27212\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27188\,
            in1 => \N__27173\,
            in2 => \N__27158\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27680\,
            in1 => \N__27665\,
            in2 => \N__27653\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27641\,
            in2 => \N__27614\,
            in3 => \N__27629\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27602\,
            in1 => \N__27587\,
            in2 => \N__27575\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27563\,
            in1 => \N__27548\,
            in2 => \N__27536\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27527\,
            in1 => \N__27512\,
            in2 => \N__27500\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27491\,
            in2 => \N__27464\,
            in3 => \N__27479\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27452\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_c_RNO_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__37976\,
            in1 => \N__37949\,
            in2 => \_gnd_net_\,
            in3 => \N__40184\,
            lcout => \current_shift_inst.un38_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_c_RNO_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40183\,
            in1 => \N__37259\,
            in2 => \_gnd_net_\,
            in3 => \N__37232\,
            lcout => \current_shift_inst.un38_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_c_RNO_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40182\,
            in1 => \N__37300\,
            in2 => \_gnd_net_\,
            in3 => \N__37274\,
            lcout => \current_shift_inst.un38_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_c_THRU_CRY_0_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40143\,
            in2 => \N__40269\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_c_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31907\,
            in2 => \N__39865\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.un38_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_c_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29150\,
            in2 => \N__40270\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0\,
            carryout => \current_shift_inst.un38_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_c_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32069\,
            in2 => \N__40219\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1\,
            carryout => \current_shift_inst.un38_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_c_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27692\,
            in2 => \N__40271\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2\,
            carryout => \current_shift_inst.un38_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_c_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27686\,
            in2 => \N__40220\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3\,
            carryout => \current_shift_inst.un38_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_c_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32144\,
            in2 => \N__40272\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4\,
            carryout => \current_shift_inst.un38_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_c_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31895\,
            in2 => \N__40221\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5\,
            carryout => \current_shift_inst.un38_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_c_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27701\,
            in2 => \N__40222\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_c_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40156\,
            in2 => \N__32126\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_7\,
            carryout => \current_shift_inst.un38_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_c_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31883\,
            in2 => \N__40223\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8\,
            carryout => \current_shift_inst.un38_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_c_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40160\,
            in2 => \N__32111\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9\,
            carryout => \current_shift_inst.un38_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_c_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37424\,
            in2 => \N__40224\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10\,
            carryout => \current_shift_inst.un38_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_c_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40164\,
            in2 => \N__32096\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11\,
            carryout => \current_shift_inst.un38_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_c_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32135\,
            in2 => \N__40225\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12\,
            carryout => \current_shift_inst.un38_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_c_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40168\,
            in2 => \N__37991\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13\,
            carryout => \current_shift_inst.un38_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_c_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32081\,
            in2 => \N__40273\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_c_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38444\,
            in2 => \N__40226\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_15\,
            carryout => \current_shift_inst.un38_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_c_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38045\,
            in2 => \N__40274\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16\,
            carryout => \current_shift_inst.un38_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_c_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40248\,
            in2 => \N__38699\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17\,
            carryout => \current_shift_inst.un38_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_c_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28622\,
            in2 => \N__40275\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18\,
            carryout => \current_shift_inst.un38_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_c_RNIBS3R1_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38759\,
            in2 => \N__40227\,
            in3 => \N__27722\,
            lcout => \current_shift_inst.control_input_1_axb_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19\,
            carryout => \current_shift_inst.un38_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_c_RNITVMS1_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38222\,
            in2 => \N__40276\,
            in3 => \N__27713\,
            lcout => \current_shift_inst.control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20\,
            carryout => \current_shift_inst.un38_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_c_RNI16PS1_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40255\,
            in2 => \N__32159\,
            in3 => \N__27704\,
            lcout => \current_shift_inst.control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21\,
            carryout => \current_shift_inst.un38_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_c_RNI5CRS1_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38852\,
            in2 => \N__40277\,
            in3 => \N__27815\,
            lcout => \current_shift_inst.control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_c_RNI9ITS1_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34127\,
            in2 => \N__40228\,
            in3 => \N__27806\,
            lcout => \current_shift_inst.control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_23\,
            carryout => \current_shift_inst.un38_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_c_RNIDOVS1_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34154\,
            in2 => \N__40278\,
            in3 => \N__27797\,
            lcout => \current_shift_inst.control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24\,
            carryout => \current_shift_inst.un38_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_c_RNIHU1T1_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34136\,
            in2 => \N__40229\,
            in3 => \N__27788\,
            lcout => \current_shift_inst.control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25\,
            carryout => \current_shift_inst.un38_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_c_RNIL44T1_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27785\,
            in2 => \N__40279\,
            in3 => \N__27767\,
            lcout => \current_shift_inst.control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26\,
            carryout => \current_shift_inst.un38_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_c_RNIPA6T1_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40265\,
            in2 => \N__32192\,
            in3 => \N__27758\,
            lcout => \current_shift_inst.control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27\,
            carryout => \current_shift_inst.un38_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_c_RNIB0AT1_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34145\,
            in2 => \N__40280\,
            in3 => \N__27749\,
            lcout => \current_shift_inst.control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28\,
            carryout => \current_shift_inst.un38_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_THRU_LUT4_0_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27746\,
            lcout => \current_shift_inst.un38_control_input_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__40181\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34007\,
            lcout => \current_shift_inst.un38_control_input_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40813\,
            in2 => \_gnd_net_\,
            in3 => \N__27929\,
            lcout => \phase_controller_inst2.time_passed_RNI9M3O\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.T01_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__27973\,
            in1 => \N__27906\,
            in2 => \_gnd_net_\,
            in3 => \N__28019\,
            lcout => \T01_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44838\,
            ce => 'H',
            sr => \N__44215\
        );

    \phase_controller_inst1.S1_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28858\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44834\,
            ce => 'H',
            sr => \N__44228\
        );

    \current_shift_inst.stop_timer_s1_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__27952\,
            in1 => \N__28857\,
            in2 => \N__28094\,
            in3 => \N__28129\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44834\,
            ce => 'H',
            sr => \N__44228\
        );

    \current_shift_inst.timer_s1.running_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__28130\,
            in1 => \N__28090\,
            in2 => \_gnd_net_\,
            in3 => \N__28112\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44834\,
            ce => 'H',
            sr => \N__44228\
        );

    \current_shift_inst.start_timer_s1_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__27951\,
            in1 => \N__28128\,
            in2 => \_gnd_net_\,
            in3 => \N__28856\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44834\,
            ce => 'H',
            sr => \N__44228\
        );

    \phase_controller_inst2.T45_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__27937\,
            in1 => \N__27844\,
            in2 => \_gnd_net_\,
            in3 => \N__27908\,
            lcout => \T45_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44834\,
            ce => 'H',
            sr => \N__44228\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28109\,
            in2 => \_gnd_net_\,
            in3 => \N__28088\,
            lcout => \current_shift_inst.timer_s1.N_166_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28110\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__28127\,
            in1 => \N__28111\,
            in2 => \_gnd_net_\,
            in3 => \N__28089\,
            lcout => \current_shift_inst.timer_s1.N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44334\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__35629\,
            in1 => \N__35828\,
            in2 => \N__32723\,
            in3 => \N__35462\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44922\,
            ce => 'H',
            sr => \N__44112\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31059\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35827\,
            in1 => \N__35630\,
            in2 => \N__35507\,
            in3 => \N__33380\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44922\,
            ce => 'H',
            sr => \N__44112\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110111"
        )
    port map (
            in0 => \N__34485\,
            in1 => \N__32245\,
            in2 => \N__32336\,
            in3 => \N__32407\,
            lcout => \current_shift_inst.PI_CTRL.N_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__28640\,
            in1 => \N__28172\,
            in2 => \N__35877\,
            in3 => \N__34283\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28208\,
            in1 => \N__28214\,
            in2 => \N__28058\,
            in3 => \N__28184\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__30287\,
            in1 => \N__28055\,
            in2 => \N__28049\,
            in3 => \N__28190\,
            lcout => \current_shift_inst.PI_CTRL.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30286\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__31241\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30630\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__30421\,
            in1 => \N__31085\,
            in2 => \N__28193\,
            in3 => \N__34645\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__34227\,
            in1 => \N__32507\,
            in2 => \_gnd_net_\,
            in3 => \N__28202\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30791\,
            in1 => \N__35321\,
            in2 => \N__34527\,
            in3 => \N__35207\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35156\,
            in1 => \N__32549\,
            in2 => \N__35042\,
            in3 => \N__34340\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__28166\,
            in1 => \N__28154\,
            in2 => \N__34172\,
            in3 => \N__28136\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__30463\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34873\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30422\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35206\,
            in1 => \N__30790\,
            in2 => \N__35328\,
            in3 => \N__34517\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34381\,
            in1 => \N__35810\,
            in2 => \N__30524\,
            in3 => \N__30893\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30685\,
            in1 => \N__30994\,
            in2 => \N__32617\,
            in3 => \N__30367\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__28519\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34877\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__34879\,
            in1 => \N__30368\,
            in2 => \N__28196\,
            in3 => \N__28505\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30686\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__30558\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34876\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30739\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__31187\,
            in1 => \N__32556\,
            in2 => \N__28478\,
            in3 => \N__34880\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30967\,
            in2 => \_gnd_net_\,
            in3 => \N__34884\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__28291\,
            in1 => \N__32251\,
            in2 => \N__34943\,
            in3 => \N__28325\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28290\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30769\,
            in2 => \_gnd_net_\,
            in3 => \N__34885\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28269\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__30928\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34883\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__34886\,
            in1 => \N__32443\,
            in2 => \N__28370\,
            in3 => \N__28270\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28238\,
            in2 => \_gnd_net_\,
            in3 => \N__28252\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28220\,
            in2 => \_gnd_net_\,
            in3 => \N__28231\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28406\,
            in2 => \_gnd_net_\,
            in3 => \N__28423\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28393\,
            in1 => \N__28382\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28376\,
            in2 => \_gnd_net_\,
            in3 => \N__28361\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28358\,
            in2 => \_gnd_net_\,
            in3 => \N__28343\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28340\,
            in2 => \_gnd_net_\,
            in3 => \N__28334\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28331\,
            in2 => \_gnd_net_\,
            in3 => \N__28319\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28316\,
            in2 => \_gnd_net_\,
            in3 => \N__28310\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_8\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28307\,
            in2 => \_gnd_net_\,
            in3 => \N__28301\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28685\,
            in2 => \_gnd_net_\,
            in3 => \N__28454\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28676\,
            in2 => \_gnd_net_\,
            in3 => \N__28451\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30464\,
            in2 => \_gnd_net_\,
            in3 => \N__28448\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31111\,
            in2 => \_gnd_net_\,
            in3 => \N__28445\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31033\,
            in2 => \_gnd_net_\,
            in3 => \N__28442\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31348\,
            in2 => \_gnd_net_\,
            in3 => \N__28439\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30559\,
            in2 => \_gnd_net_\,
            in3 => \N__28436\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30929\,
            in2 => \_gnd_net_\,
            in3 => \N__28433\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30847\,
            in2 => \_gnd_net_\,
            in3 => \N__28430\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28520\,
            in2 => \_gnd_net_\,
            in3 => \N__28496\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30770\,
            in2 => \_gnd_net_\,
            in3 => \N__28493\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30968\,
            in2 => \_gnd_net_\,
            in3 => \N__28490\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31936\,
            in2 => \_gnd_net_\,
            in3 => \N__28487\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30740\,
            in2 => \_gnd_net_\,
            in3 => \N__28484\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31293\,
            in2 => \_gnd_net_\,
            in3 => \N__28481\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31186\,
            in2 => \_gnd_net_\,
            in3 => \N__28463\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30595\,
            in3 => \N__28460\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33264\,
            in2 => \_gnd_net_\,
            in3 => \N__28457\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31137\,
            in2 => \_gnd_net_\,
            in3 => \N__28610\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33516\,
            in2 => \_gnd_net_\,
            in3 => \N__28607\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31957\,
            in2 => \_gnd_net_\,
            in3 => \N__28604\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__34833\,
            in1 => \N__28663\,
            in2 => \_gnd_net_\,
            in3 => \N__28601\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIL7IU_0_1_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__28553\,
            in1 => \N__44318\,
            in2 => \N__28597\,
            in3 => \N__43178\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__43179\,
            in1 => \N__28596\,
            in2 => \N__43143\,
            in3 => \N__28554\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44876\,
            ce => 'H',
            sr => \N__44150\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43174\,
            in2 => \_gnd_net_\,
            in3 => \N__43132\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001100100"
        )
    port map (
            in0 => \N__28555\,
            in1 => \N__43181\,
            in2 => \N__28598\,
            in3 => \N__43139\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44876\,
            ce => 'H',
            sr => \N__44150\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIL7IU_1_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101110"
        )
    port map (
            in0 => \N__44319\,
            in1 => \N__28589\,
            in2 => \N__43188\,
            in3 => \N__28552\,
            lcout => \phase_controller_inst1.stoper_tr.un1_stoper_state12_1_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000010"
        )
    port map (
            in0 => \N__43180\,
            in1 => \N__28532\,
            in2 => \N__43144\,
            in3 => \N__28725\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44876\,
            ce => 'H',
            sr => \N__44150\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__31462\,
            in1 => \N__28705\,
            in2 => \_gnd_net_\,
            in3 => \N__28808\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44869\,
            ce => 'H',
            sr => \N__31407\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34993\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30249\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35878\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30908\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28662\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34584\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_c_RNO_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40115\,
            in1 => \_gnd_net_\,
            in2 => \N__38123\,
            in3 => \N__38093\,
            lcout => \current_shift_inst.un38_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38118\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_c_RNO_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__40114\,
            in1 => \N__33755\,
            in2 => \_gnd_net_\,
            in3 => \N__33806\,
            lcout => \current_shift_inst.un38_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__29055\,
            in1 => \N__29144\,
            in2 => \_gnd_net_\,
            in3 => \N__29108\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44863\,
            ce => 'H',
            sr => \N__44160\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29054\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__36017\,
            in1 => \N__36553\,
            in2 => \N__37180\,
            in3 => \N__36182\,
            lcout => \elapsed_time_ns_1_RNIAE2591_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_2_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__28894\,
            in1 => \N__36588\,
            in2 => \N__36632\,
            in3 => \N__28859\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44858\,
            ce => 'H',
            sr => \N__44169\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_0_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__32023\,
            in1 => \N__32050\,
            in2 => \N__28813\,
            in3 => \N__31457\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44858\,
            ce => 'H',
            sr => \N__44169\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_1_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001000000010"
        )
    port map (
            in0 => \N__31456\,
            in1 => \N__28804\,
            in2 => \N__32057\,
            in3 => \N__32024\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44858\,
            ce => 'H',
            sr => \N__44169\
        );

    \phase_controller_inst1.state_1_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__29403\,
            in1 => \N__36589\,
            in2 => \N__28769\,
            in3 => \N__36630\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44858\,
            ce => 'H',
            sr => \N__44169\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29368\,
            in2 => \N__33649\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__44854\,
            ce => \N__38178\,
            sr => \N__44177\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29343\,
            in2 => \N__33841\,
            in3 => \N__29177\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__44854\,
            ce => \N__38178\,
            sr => \N__44177\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29369\,
            in2 => \N__29321\,
            in3 => \N__29174\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__44854\,
            ce => \N__38178\,
            sr => \N__44177\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29287\,
            in2 => \N__29348\,
            in3 => \N__29171\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__44854\,
            ce => \N__38178\,
            sr => \N__44177\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29320\,
            in2 => \N__29260\,
            in3 => \N__29168\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__44854\,
            ce => \N__38178\,
            sr => \N__44177\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29644\,
            in2 => \N__29291\,
            in3 => \N__29165\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__44854\,
            ce => \N__38178\,
            sr => \N__44177\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29614\,
            in2 => \N__29261\,
            in3 => \N__29162\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__44854\,
            ce => \N__38178\,
            sr => \N__44177\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29645\,
            in2 => \N__29584\,
            in3 => \N__29159\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__44854\,
            ce => \N__38178\,
            sr => \N__44177\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29551\,
            in2 => \N__29621\,
            in3 => \N__29156\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__44850\,
            ce => \N__38177\,
            sr => \N__44180\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29527\,
            in2 => \N__29588\,
            in3 => \N__29153\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__44850\,
            ce => \N__38177\,
            sr => \N__44180\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29552\,
            in2 => \N__29506\,
            in3 => \N__29204\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__44850\,
            ce => \N__38177\,
            sr => \N__44180\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29528\,
            in2 => \N__29476\,
            in3 => \N__29201\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__44850\,
            ce => \N__38177\,
            sr => \N__44180\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29443\,
            in2 => \N__29507\,
            in3 => \N__29198\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__44850\,
            ce => \N__38177\,
            sr => \N__44180\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29899\,
            in2 => \N__29477\,
            in3 => \N__29195\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__44850\,
            ce => \N__38177\,
            sr => \N__44180\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29872\,
            in2 => \N__29447\,
            in3 => \N__29192\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__44850\,
            ce => \N__38177\,
            sr => \N__44180\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29900\,
            in2 => \N__29842\,
            in3 => \N__29189\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__44850\,
            ce => \N__38177\,
            sr => \N__44180\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29806\,
            in2 => \N__29876\,
            in3 => \N__29186\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__44847\,
            ce => \N__38176\,
            sr => \N__44187\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29782\,
            in2 => \N__29843\,
            in3 => \N__29183\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__44847\,
            ce => \N__38176\,
            sr => \N__44187\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29807\,
            in2 => \N__29761\,
            in3 => \N__29180\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__44847\,
            ce => \N__38176\,
            sr => \N__44187\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29783\,
            in2 => \N__29731\,
            in3 => \N__29231\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__44847\,
            ce => \N__38176\,
            sr => \N__44187\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29698\,
            in2 => \N__29762\,
            in3 => \N__29228\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__44847\,
            ce => \N__38176\,
            sr => \N__44187\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29671\,
            in2 => \N__29732\,
            in3 => \N__29225\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__44847\,
            ce => \N__38176\,
            sr => \N__44187\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30202\,
            in2 => \N__29702\,
            in3 => \N__29222\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__44847\,
            ce => \N__38176\,
            sr => \N__44187\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30175\,
            in2 => \N__29675\,
            in3 => \N__29219\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__44847\,
            ce => \N__38176\,
            sr => \N__44187\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30148\,
            in2 => \N__30206\,
            in3 => \N__29216\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_13_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__44844\,
            ce => \N__38175\,
            sr => \N__44201\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30124\,
            in2 => \N__30179\,
            in3 => \N__29213\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__44844\,
            ce => \N__38175\,
            sr => \N__44201\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30149\,
            in2 => \N__30104\,
            in3 => \N__29210\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__44844\,
            ce => \N__38175\,
            sr => \N__44201\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30125\,
            in2 => \N__29957\,
            in3 => \N__29207\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__44844\,
            ce => \N__38175\,
            sr => \N__44201\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29417\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29412\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44842\,
            ce => 'H',
            sr => \N__44209\
        );

    \current_shift_inst.timer_s1.counter_0_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30073\,
            in1 => \N__33633\,
            in2 => \_gnd_net_\,
            in3 => \N__29375\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__44840\,
            ce => \N__29936\,
            sr => \N__44216\
        );

    \current_shift_inst.timer_s1.counter_1_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30069\,
            in1 => \N__33825\,
            in2 => \_gnd_net_\,
            in3 => \N__29372\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__44840\,
            ce => \N__29936\,
            sr => \N__44216\
        );

    \current_shift_inst.timer_s1.counter_2_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30074\,
            in1 => \N__29367\,
            in2 => \_gnd_net_\,
            in3 => \N__29351\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__44840\,
            ce => \N__29936\,
            sr => \N__44216\
        );

    \current_shift_inst.timer_s1.counter_3_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30070\,
            in1 => \N__29347\,
            in2 => \_gnd_net_\,
            in3 => \N__29324\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__44840\,
            ce => \N__29936\,
            sr => \N__44216\
        );

    \current_shift_inst.timer_s1.counter_4_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30075\,
            in1 => \N__29310\,
            in2 => \_gnd_net_\,
            in3 => \N__29294\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__44840\,
            ce => \N__29936\,
            sr => \N__44216\
        );

    \current_shift_inst.timer_s1.counter_5_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30071\,
            in1 => \N__29280\,
            in2 => \_gnd_net_\,
            in3 => \N__29264\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__44840\,
            ce => \N__29936\,
            sr => \N__44216\
        );

    \current_shift_inst.timer_s1.counter_6_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30076\,
            in1 => \N__29248\,
            in2 => \_gnd_net_\,
            in3 => \N__29234\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__44840\,
            ce => \N__29936\,
            sr => \N__44216\
        );

    \current_shift_inst.timer_s1.counter_7_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30072\,
            in1 => \N__29638\,
            in2 => \_gnd_net_\,
            in3 => \N__29624\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__44840\,
            ce => \N__29936\,
            sr => \N__44216\
        );

    \current_shift_inst.timer_s1.counter_8_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30049\,
            in1 => \N__29613\,
            in2 => \_gnd_net_\,
            in3 => \N__29591\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__44837\,
            ce => \N__29931\,
            sr => \N__44223\
        );

    \current_shift_inst.timer_s1.counter_9_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30053\,
            in1 => \N__29577\,
            in2 => \_gnd_net_\,
            in3 => \N__29555\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__44837\,
            ce => \N__29931\,
            sr => \N__44223\
        );

    \current_shift_inst.timer_s1.counter_10_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30046\,
            in1 => \N__29545\,
            in2 => \_gnd_net_\,
            in3 => \N__29531\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__44837\,
            ce => \N__29931\,
            sr => \N__44223\
        );

    \current_shift_inst.timer_s1.counter_11_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30050\,
            in1 => \N__29526\,
            in2 => \_gnd_net_\,
            in3 => \N__29510\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__44837\,
            ce => \N__29931\,
            sr => \N__44223\
        );

    \current_shift_inst.timer_s1.counter_12_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30047\,
            in1 => \N__29494\,
            in2 => \_gnd_net_\,
            in3 => \N__29480\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__44837\,
            ce => \N__29931\,
            sr => \N__44223\
        );

    \current_shift_inst.timer_s1.counter_13_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30051\,
            in1 => \N__29464\,
            in2 => \_gnd_net_\,
            in3 => \N__29450\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__44837\,
            ce => \N__29931\,
            sr => \N__44223\
        );

    \current_shift_inst.timer_s1.counter_14_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30048\,
            in1 => \N__29436\,
            in2 => \_gnd_net_\,
            in3 => \N__29420\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__44837\,
            ce => \N__29931\,
            sr => \N__44223\
        );

    \current_shift_inst.timer_s1.counter_15_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30052\,
            in1 => \N__29893\,
            in2 => \_gnd_net_\,
            in3 => \N__29879\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__44837\,
            ce => \N__29931\,
            sr => \N__44223\
        );

    \current_shift_inst.timer_s1.counter_16_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30077\,
            in1 => \N__29865\,
            in2 => \_gnd_net_\,
            in3 => \N__29846\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__44835\,
            ce => \N__29930\,
            sr => \N__44229\
        );

    \current_shift_inst.timer_s1.counter_17_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30042\,
            in1 => \N__29829\,
            in2 => \_gnd_net_\,
            in3 => \N__29810\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__44835\,
            ce => \N__29930\,
            sr => \N__44229\
        );

    \current_shift_inst.timer_s1.counter_18_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30078\,
            in1 => \N__29800\,
            in2 => \_gnd_net_\,
            in3 => \N__29786\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__44835\,
            ce => \N__29930\,
            sr => \N__44229\
        );

    \current_shift_inst.timer_s1.counter_19_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30043\,
            in1 => \N__29781\,
            in2 => \_gnd_net_\,
            in3 => \N__29765\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__44835\,
            ce => \N__29930\,
            sr => \N__44229\
        );

    \current_shift_inst.timer_s1.counter_20_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30079\,
            in1 => \N__29749\,
            in2 => \_gnd_net_\,
            in3 => \N__29735\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__44835\,
            ce => \N__29930\,
            sr => \N__44229\
        );

    \current_shift_inst.timer_s1.counter_21_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30044\,
            in1 => \N__29719\,
            in2 => \_gnd_net_\,
            in3 => \N__29705\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__44835\,
            ce => \N__29930\,
            sr => \N__44229\
        );

    \current_shift_inst.timer_s1.counter_22_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30080\,
            in1 => \N__29697\,
            in2 => \_gnd_net_\,
            in3 => \N__29678\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__44835\,
            ce => \N__29930\,
            sr => \N__44229\
        );

    \current_shift_inst.timer_s1.counter_23_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30045\,
            in1 => \N__29664\,
            in2 => \_gnd_net_\,
            in3 => \N__29648\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__44835\,
            ce => \N__29930\,
            sr => \N__44229\
        );

    \current_shift_inst.timer_s1.counter_24_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30054\,
            in1 => \N__30201\,
            in2 => \_gnd_net_\,
            in3 => \N__30182\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_13_27_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__44832\,
            ce => \N__29932\,
            sr => \N__44232\
        );

    \current_shift_inst.timer_s1.counter_25_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30058\,
            in1 => \N__30168\,
            in2 => \_gnd_net_\,
            in3 => \N__30152\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__44832\,
            ce => \N__29932\,
            sr => \N__44232\
        );

    \current_shift_inst.timer_s1.counter_26_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30055\,
            in1 => \N__30142\,
            in2 => \_gnd_net_\,
            in3 => \N__30128\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__44832\,
            ce => \N__29932\,
            sr => \N__44232\
        );

    \current_shift_inst.timer_s1.counter_27_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30059\,
            in1 => \N__30123\,
            in2 => \_gnd_net_\,
            in3 => \N__30107\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__44832\,
            ce => \N__29932\,
            sr => \N__44232\
        );

    \current_shift_inst.timer_s1.counter_28_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30056\,
            in1 => \N__30097\,
            in2 => \_gnd_net_\,
            in3 => \N__30083\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__44832\,
            ce => \N__29932\,
            sr => \N__44232\
        );

    \current_shift_inst.timer_s1.counter_29_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__29950\,
            in1 => \N__30057\,
            in2 => \_gnd_net_\,
            in3 => \N__29960\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44832\,
            ce => \N__29932\,
            sr => \N__44232\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32533\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32491\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000111110101"
        )
    port map (
            in0 => \N__35826\,
            in1 => \N__35632\,
            in2 => \N__35509\,
            in3 => \N__32681\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44929\,
            ce => 'H',
            sr => \N__44107\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000111110101"
        )
    port map (
            in0 => \N__35825\,
            in1 => \N__35631\,
            in2 => \N__35508\,
            in3 => \N__32780\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44929\,
            ce => 'H',
            sr => \N__44107\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__30294\,
            in1 => \N__34947\,
            in2 => \N__30344\,
            in3 => \N__30314\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35588\,
            in1 => \N__35832\,
            in2 => \N__32822\,
            in3 => \N__35445\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44923\,
            ce => 'H',
            sr => \N__44113\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35829\,
            in1 => \N__35589\,
            in2 => \N__35494\,
            in3 => \N__33017\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44923\,
            ce => 'H',
            sr => \N__44113\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35586\,
            in1 => \N__35830\,
            in2 => \N__32987\,
            in3 => \N__35443\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44923\,
            ce => 'H',
            sr => \N__44113\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35587\,
            in1 => \N__35831\,
            in2 => \N__32966\,
            in3 => \N__35444\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44923\,
            ce => 'H',
            sr => \N__44113\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34386\,
            in1 => \N__35867\,
            in2 => \N__30523\,
            in3 => \N__30892\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__30626\,
            in1 => \N__30251\,
            in2 => \N__34964\,
            in3 => \N__30218\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30625\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001110101111"
        )
    port map (
            in0 => \N__35431\,
            in1 => \N__35635\,
            in2 => \N__35833\,
            in3 => \N__32753\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44917\,
            ce => 'H',
            sr => \N__44117\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__32936\,
            in1 => \N__35813\,
            in2 => \N__35672\,
            in3 => \N__35432\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44917\,
            ce => 'H',
            sr => \N__44117\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35811\,
            in1 => \N__35633\,
            in2 => \N__35492\,
            in3 => \N__32906\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44917\,
            ce => 'H',
            sr => \N__44117\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__32876\,
            in1 => \N__35814\,
            in2 => \N__35671\,
            in3 => \N__35439\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44917\,
            ce => 'H',
            sr => \N__44117\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35812\,
            in1 => \N__35634\,
            in2 => \N__35493\,
            in3 => \N__32849\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44917\,
            ce => 'H',
            sr => \N__44117\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__30602\,
            in1 => \N__32509\,
            in2 => \N__34961\,
            in3 => \N__30572\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__30560\,
            in1 => \N__30528\,
            in2 => \N__30479\,
            in3 => \N__34933\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__30462\,
            in1 => \N__30439\,
            in2 => \N__34959\,
            in3 => \N__30392\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30369\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011111111"
        )
    port map (
            in0 => \N__30995\,
            in1 => \N__30966\,
            in2 => \N__30947\,
            in3 => \N__34938\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__30927\,
            in1 => \N__30900\,
            in2 => \N__34960\,
            in3 => \N__30863\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__34390\,
            in1 => \N__34937\,
            in2 => \N__30851\,
            in3 => \N__30821\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__30804\,
            in1 => \N__30768\,
            in2 => \N__34954\,
            in3 => \N__30749\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32406\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35043\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__34341\,
            in1 => \N__30738\,
            in2 => \N__34955\,
            in3 => \N__30719\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__31937\,
            in1 => \N__30702\,
            in2 => \N__30662\,
            in3 => \N__34926\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__31267\,
            in1 => \N__31225\,
            in2 => \N__34953\,
            in3 => \N__31196\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35217\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34899\,
            in2 => \_gnd_net_\,
            in3 => \N__31185\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__31961\,
            in1 => \N__35047\,
            in2 => \N__34949\,
            in3 => \N__31160\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__35170\,
            in1 => \N__34905\,
            in2 => \N__31148\,
            in3 => \N__31121\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34897\,
            in1 => \N__31112\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__31095\,
            in1 => \N__34901\,
            in2 => \N__31043\,
            in3 => \N__31040\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34898\,
            in1 => \N__31034\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__35329\,
            in1 => \N__34900\,
            in2 => \N__31022\,
            in3 => \N__31019\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__31349\,
            in1 => \N__34222\,
            in2 => \N__34948\,
            in3 => \N__31319\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100100"
        )
    port map (
            in0 => \N__36513\,
            in1 => \N__42488\,
            in2 => \N__39245\,
            in3 => \N__36363\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__36309\,
            in1 => \_gnd_net_\,
            in2 => \N__31313\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIFG4DM1_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__36509\,
            in1 => \N__39368\,
            in2 => \N__33467\,
            in3 => \N__36152\,
            lcout => \elapsed_time_ns_1_RNIRBJF91_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111101010"
        )
    port map (
            in0 => \N__36308\,
            in1 => \N__36512\,
            in2 => \N__38660\,
            in3 => \N__37078\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31310\,
            in3 => \N__36362\,
            lcout => \elapsed_time_ns_1_RNIRHL2M1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__34872\,
            in1 => \N__32608\,
            in2 => \N__31307\,
            in3 => \N__31280\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__36511\,
            in1 => \N__38954\,
            in2 => \N__42535\,
            in3 => \N__36153\,
            lcout => \elapsed_time_ns_1_RNIQ8HF91_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__39134\,
            in1 => \N__36510\,
            in2 => \N__36172\,
            in3 => \N__33440\,
            lcout => \elapsed_time_ns_1_RNIQ9IF91_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__38975\,
            in1 => \N__36516\,
            in2 => \N__36177\,
            in3 => \N__41517\,
            lcout => \elapsed_time_ns_1_RNIP7HF91_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__36041\,
            in1 => \N__44313\,
            in2 => \_gnd_net_\,
            in3 => \N__33551\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__44314\,
            in1 => \N__39338\,
            in2 => \N__31364\,
            in3 => \N__33557\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31361\,
            in3 => \N__31355\,
            lcout => \elapsed_time_ns_1_RNIHI4DM1_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__36922\,
            in1 => \N__36517\,
            in2 => \N__39011\,
            in3 => \N__36385\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31358\,
            in3 => \N__36310\,
            lcout => \elapsed_time_ns_1_RNI1OL2M1_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__33287\,
            in1 => \_gnd_net_\,
            in2 => \N__36321\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIUKL2M1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__36518\,
            in1 => \N__39188\,
            in2 => \N__36396\,
            in3 => \N__42330\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33563\,
            in2 => \_gnd_net_\,
            in3 => \N__36314\,
            lcout => \elapsed_time_ns_1_RNIIJ4DM1_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__39068\,
            in1 => \N__36167\,
            in2 => \N__36867\,
            in3 => \N__36524\,
            lcout => \elapsed_time_ns_1_RNIFJ2591_0_7\,
            ltout => \elapsed_time_ns_1_RNIFJ2591_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_2_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__36794\,
            in1 => \N__36836\,
            in2 => \N__31871\,
            in3 => \N__36898\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_6_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__42006\,
            in1 => \_gnd_net_\,
            in2 => \N__31868\,
            in3 => \N__37020\,
            lcout => \phase_controller_inst1.stoper_tr.N_250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__31865\,
            in1 => \N__31691\,
            in2 => \N__31657\,
            in3 => \N__31577\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_0_a5_1_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__42007\,
            in1 => \N__37112\,
            in2 => \N__37154\,
            in3 => \N__31970\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.N_235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_0_1_1_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33690\,
            in2 => \N__31535\,
            in3 => \N__36751\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_f0_0_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0_3_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__42069\,
            in1 => \N__42167\,
            in2 => \N__37120\,
            in3 => \N__37146\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_3_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__37086\,
            in1 => \N__37619\,
            in2 => \N__31532\,
            in3 => \N__36770\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44883\,
            ce => \N__43743\,
            sr => \N__44144\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_RNI74R51_0_1_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__32056\,
            in1 => \N__44316\,
            in2 => \N__31471\,
            in3 => \N__32029\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_RNI74R51_1_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111110"
        )
    port map (
            in0 => \N__44317\,
            in1 => \N__32055\,
            in2 => \N__32030\,
            in3 => \N__31463\,
            lcout => \phase_controller_inst2.stoper_hc.un1_stoper_state12_1_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32054\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32025\,
            lcout => \phase_controller_inst2.stoper_hc.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_0_o2_1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__37079\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37170\,
            lcout => \phase_controller_inst1.stoper_tr.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34916\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31956\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31929\,
            in2 => \_gnd_net_\,
            in3 => \N__34915\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32613\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33612\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_c_RNO_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100011101"
        )
    port map (
            in0 => \N__33613\,
            in1 => \N__40061\,
            in2 => \N__31910\,
            in3 => \N__39857\,
            lcout => \current_shift_inst.un38_control_input_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_c_RNO_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40117\,
            in1 => \N__37376\,
            in2 => \_gnd_net_\,
            in3 => \N__37352\,
            lcout => \current_shift_inst.un38_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_c_RNO_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__37934\,
            in1 => \N__40119\,
            in2 => \_gnd_net_\,
            in3 => \N__37904\,
            lcout => \current_shift_inst.un38_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_c_RNO_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40118\,
            in1 => \_gnd_net_\,
            in2 => \N__37339\,
            in3 => \N__37313\,
            lcout => \current_shift_inst.un38_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_c_RNO_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__37660\,
            in1 => \N__40120\,
            in2 => \_gnd_net_\,
            in3 => \N__37634\,
            lcout => \current_shift_inst.un38_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_c_RNO_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40121\,
            in1 => \N__37891\,
            in2 => \_gnd_net_\,
            in3 => \N__37865\,
            lcout => \current_shift_inst.un38_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_c_RNO_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__37835\,
            in1 => \N__40122\,
            in2 => \_gnd_net_\,
            in3 => \N__37847\,
            lcout => \current_shift_inst.un38_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_c_RNO_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40116\,
            in1 => \N__37400\,
            in2 => \_gnd_net_\,
            in3 => \N__37412\,
            lcout => \current_shift_inst.un38_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37332\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37449\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37920\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37387\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37363\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40124\,
            in1 => \N__38263\,
            in2 => \_gnd_net_\,
            in3 => \N__38236\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37290\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37245\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_c_RNO_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__37450\,
            in1 => \N__40123\,
            in2 => \_gnd_net_\,
            in3 => \N__37436\,
            lcout => \current_shift_inst.un38_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_c_RNO_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40057\,
            in1 => \N__37762\,
            in2 => \_gnd_net_\,
            in3 => \N__37742\,
            lcout => \current_shift_inst.un38_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__37730\,
            in1 => \N__38473\,
            in2 => \_gnd_net_\,
            in3 => \N__38455\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37650\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38017\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37881\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38472\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37794\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38739\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__43838\,
            in1 => \N__44378\,
            in2 => \_gnd_net_\,
            in3 => \N__43671\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44855\,
            ce => 'H',
            sr => \N__44588\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37962\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38143\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37758\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38056\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_1_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__33698\,
            in1 => \N__37620\,
            in2 => \N__42267\,
            in3 => \N__33671\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44851\,
            ce => \N__41941\,
            sr => \N__44181\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_4_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__37622\,
            in1 => \N__42252\,
            in2 => \N__37502\,
            in3 => \N__37540\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44851\,
            ce => \N__41941\,
            sr => \N__44181\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_3_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__32168\,
            in1 => \N__37621\,
            in2 => \N__36775\,
            in3 => \N__37091\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44851\,
            ce => \N__41941\,
            sr => \N__44181\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__40063\,
            in1 => \_gnd_net_\,
            in2 => \N__34037\,
            in3 => \N__32180\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32179\,
            in1 => \N__40062\,
            in2 => \_gnd_net_\,
            in3 => \N__34033\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32178\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38295\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38830\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38536\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38373\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38418\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35818\,
            in1 => \N__35644\,
            in2 => \N__35510\,
            in3 => \N__33227\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44934\,
            ce => 'H',
            sr => \N__44105\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35642\,
            in1 => \N__35820\,
            in2 => \N__33188\,
            in3 => \N__35475\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44934\,
            ce => 'H',
            sr => \N__44105\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35819\,
            in1 => \N__35645\,
            in2 => \N__35511\,
            in3 => \N__33146\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44934\,
            ce => 'H',
            sr => \N__44105\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35643\,
            in1 => \N__35821\,
            in2 => \N__33113\,
            in3 => \N__35476\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44934\,
            ce => 'H',
            sr => \N__44105\
        );

    \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32461\,
            in2 => \N__32465\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__35675\,
            in1 => \N__32444\,
            in2 => \N__32429\,
            in3 => \N__32375\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            clk => \N__44930\,
            ce => 'H',
            sr => \N__44108\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__35677\,
            in1 => \N__32372\,
            in2 => \N__32360\,
            in3 => \N__32300\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            clk => \N__44930\,
            ce => 'H',
            sr => \N__44108\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__35676\,
            in1 => \N__32297\,
            in2 => \N__34409\,
            in3 => \N__32285\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            clk => \N__44930\,
            ce => 'H',
            sr => \N__44108\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0111110111010111"
        )
    port map (
            in0 => \N__35678\,
            in1 => \N__32282\,
            in2 => \N__32270\,
            in3 => \N__32204\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            clk => \N__44930\,
            ce => 'H',
            sr => \N__44108\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32201\,
            in2 => \N__32834\,
            in3 => \N__32810\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32807\,
            in2 => \N__32795\,
            in3 => \N__32774\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34265\,
            in2 => \N__34670\,
            in3 => \N__32771\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32768\,
            in2 => \N__32762\,
            in3 => \N__32744\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32741\,
            in2 => \N__32732\,
            in3 => \N__32708\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32705\,
            in2 => \N__32696\,
            in3 => \N__32672\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34259\,
            in2 => \N__32669\,
            in3 => \N__32654\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32651\,
            in2 => \N__32636\,
            in3 => \N__32621\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33038\,
            in2 => \N__33026\,
            in3 => \N__33011\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33008\,
            in2 => \N__32996\,
            in3 => \N__32978\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34352\,
            in2 => \N__32975\,
            in3 => \N__32957\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32954\,
            in2 => \N__32948\,
            in3 => \N__32930\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32927\,
            in2 => \N__32915\,
            in3 => \N__32900\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32897\,
            in2 => \N__32885\,
            in3 => \N__32870\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32867\,
            in2 => \N__32858\,
            in3 => \N__32843\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32840\,
            in2 => \N__34295\,
            in3 => \N__33218\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33215\,
            in2 => \N__33200\,
            in3 => \N__33176\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33173\,
            in2 => \N__33161\,
            in3 => \N__33137\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33134\,
            in2 => \N__33122\,
            in3 => \N__33098\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33233\,
            in2 => \N__33095\,
            in3 => \N__33086\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34274\,
            in2 => \N__33083\,
            in3 => \N__33074\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33071\,
            in2 => \N__33491\,
            in3 => \N__33059\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33056\,
            in2 => \N__33050\,
            in3 => \N__33041\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33413\,
            in2 => \N__33398\,
            in3 => \N__33368\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33330\,
            in2 => \N__33365\,
            in3 => \N__33350\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33332\,
            in2 => \N__33347\,
            in3 => \N__33335\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33331\,
            in2 => \N__33311\,
            in3 => \N__33293\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__34914\,
            in1 => \N__35778\,
            in2 => \_gnd_net_\,
            in3 => \N__33290\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__36815\,
            in1 => \N__36530\,
            in2 => \N__38582\,
            in3 => \N__36370\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__39268\,
            in1 => \N__35243\,
            in2 => \N__38887\,
            in3 => \N__35996\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__39342\,
            in1 => \N__36249\,
            in2 => \N__33278\,
            in3 => \N__36266\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011111111"
        )
    port map (
            in0 => \N__35221\,
            in1 => \N__33275\,
            in2 => \N__33248\,
            in3 => \N__34912\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__35110\,
            in1 => \N__34913\,
            in2 => \N__33530\,
            in3 => \N__33503\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__36145\,
            in1 => \N__33452\,
            in2 => \N__39116\,
            in3 => \N__36507\,
            lcout => \elapsed_time_ns_1_RNIRAIF91_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__35914\,
            in1 => \N__44311\,
            in2 => \N__36376\,
            in3 => \N__35273\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__44312\,
            in1 => \N__39344\,
            in2 => \N__33479\,
            in3 => \N__36040\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\,
            ltout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__36508\,
            in1 => \N__38933\,
            in2 => \N__33476\,
            in3 => \N__41592\,
            lcout => \elapsed_time_ns_1_RNIR9HF91_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__33428\,
            in1 => \N__36506\,
            in2 => \N__36171\,
            in3 => \N__39092\,
            lcout => \elapsed_time_ns_1_RNISBIF91_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__39392\,
            in1 => \N__33473\,
            in2 => \N__36543\,
            in3 => \N__36144\,
            lcout => \elapsed_time_ns_1_RNI3JIF91_0_29\,
            ltout => \elapsed_time_ns_1_RNI3JIF91_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_o5_7_15_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33463\,
            in1 => \N__33451\,
            in2 => \N__33443\,
            in3 => \N__33439\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_7_i_o5_7Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_o5_15_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35981\,
            in1 => \N__33427\,
            in2 => \N__33416\,
            in3 => \N__36203\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__35920\,
            in1 => \N__36250\,
            in2 => \N__35960\,
            in3 => \N__36264\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_359_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__36156\,
            in1 => \N__36520\,
            in2 => \N__39044\,
            in3 => \N__36841\,
            lcout => \elapsed_time_ns_1_RNIGK2591_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__35272\,
            in1 => \N__36251\,
            in2 => \N__35924\,
            in3 => \N__36265\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_381\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__36036\,
            in1 => \N__33550\,
            in2 => \N__33539\,
            in3 => \N__39337\,
            lcout => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\,
            ltout => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__38912\,
            in1 => \N__42396\,
            in2 => \N__33536\,
            in3 => \N__36154\,
            lcout => \elapsed_time_ns_1_RNISAHF91_0_13\,
            ltout => \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_a2_2_2_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41585\,
            in1 => \N__41511\,
            in2 => \N__33533\,
            in3 => \N__42521\,
            lcout => \phase_controller_inst1.stoper_tr.N_244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__36307\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33572\,
            lcout => \elapsed_time_ns_1_RNIGH4DM1_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__36155\,
            in1 => \N__36519\,
            in2 => \N__37539\,
            in3 => \N__38627\,
            lcout => \elapsed_time_ns_1_RNICG2591_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_9_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__42324\,
            in1 => \N__42498\,
            in2 => \N__42372\,
            in3 => \N__42290\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__36515\,
            in1 => \N__36163\,
            in2 => \N__37029\,
            in3 => \N__39272\,
            lcout => \elapsed_time_ns_1_RNIUCHF91_0_15\,
            ltout => \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_9_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36917\,
            in2 => \N__33590\,
            in3 => \N__41552\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.N_251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_2_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__42499\,
            in1 => \N__42365\,
            in2 => \N__33587\,
            in3 => \N__33581\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__38606\,
            in1 => \N__36942\,
            in2 => \N__36176\,
            in3 => \N__36514\,
            lcout => \elapsed_time_ns_1_RNIDH2591_0_5\,
            ltout => \elapsed_time_ns_1_RNIDH2591_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3_2_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42289\,
            in1 => \N__42323\,
            in2 => \N__33584\,
            in3 => \N__37523\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_a2_10_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__37021\,
            in1 => \N__36968\,
            in2 => \_gnd_net_\,
            in3 => \N__41553\,
            lcout => \phase_controller_inst1.stoper_tr.N_241\,
            ltout => \phase_controller_inst1.stoper_tr.N_241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_i_1_9_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__36918\,
            in1 => \_gnd_net_\,
            in2 => \N__33575\,
            in3 => \N__42009\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__42303\,
            in1 => \N__36541\,
            in2 => \N__36397\,
            in3 => \N__39212\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__42371\,
            in1 => \N__36542\,
            in2 => \N__36398\,
            in3 => \N__39161\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001110"
        )
    port map (
            in0 => \N__36540\,
            in1 => \N__33691\,
            in2 => \N__38684\,
            in3 => \N__36389\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33701\,
            in3 => \N__36322\,
            lcout => \elapsed_time_ns_1_RNIPFL2M1_0_1\,
            ltout => \elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_1_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__42166\,
            in1 => \N__37592\,
            in2 => \N__33674\,
            in3 => \N__33664\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44889\,
            ce => \N__43736\,
            sr => \N__44138\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__39343\,
            in1 => \N__42165\,
            in2 => \N__36178\,
            in3 => \N__36539\,
            lcout => \elapsed_time_ns_1_RNISCJF91_0_31\,
            ltout => \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_a2_2_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__37022\,
            in1 => \N__37113\,
            in2 => \N__33653\,
            in3 => \N__42008\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33650\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44884\,
            ce => \N__38180\,
            sr => \N__44145\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__37693\,
            in1 => \N__33614\,
            in2 => \_gnd_net_\,
            in3 => \N__33777\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__40461\,
            in1 => \_gnd_net_\,
            in2 => \N__33599\,
            in3 => \N__33596\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__38210\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44884\,
            ce => \N__38180\,
            sr => \N__44145\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38209\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44884\,
            ce => \N__38180\,
            sr => \N__44145\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__37694\,
            in1 => \_gnd_net_\,
            in2 => \N__33754\,
            in3 => \N__33799\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33842\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44884\,
            ce => \N__38180\,
            sr => \N__44145\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33798\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33785\,
            in2 => \N__33778\,
            in3 => \N__33779\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33737\,
            in2 => \_gnd_net_\,
            in3 => \N__33731\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33728\,
            in2 => \_gnd_net_\,
            in3 => \N__33722\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33719\,
            in2 => \_gnd_net_\,
            in3 => \N__33713\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33710\,
            in2 => \_gnd_net_\,
            in3 => \N__33704\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33929\,
            in2 => \_gnd_net_\,
            in3 => \N__33923\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33920\,
            in2 => \_gnd_net_\,
            in3 => \N__33911\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33908\,
            in2 => \_gnd_net_\,
            in3 => \N__33902\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33899\,
            in2 => \_gnd_net_\,
            in3 => \N__33893\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33890\,
            in2 => \_gnd_net_\,
            in3 => \N__33884\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33881\,
            in2 => \_gnd_net_\,
            in3 => \N__33875\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33872\,
            in2 => \_gnd_net_\,
            in3 => \N__33866\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33863\,
            in2 => \_gnd_net_\,
            in3 => \N__33854\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33851\,
            in2 => \_gnd_net_\,
            in3 => \N__33845\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37853\,
            in2 => \_gnd_net_\,
            in3 => \N__33992\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33989\,
            in2 => \_gnd_net_\,
            in3 => \N__33983\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33980\,
            in2 => \_gnd_net_\,
            in3 => \N__33974\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33971\,
            in3 => \N__33962\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33959\,
            in2 => \_gnd_net_\,
            in3 => \N__33947\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34160\,
            in2 => \_gnd_net_\,
            in3 => \N__33944\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33941\,
            in2 => \_gnd_net_\,
            in3 => \N__33935\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34118\,
            in2 => \_gnd_net_\,
            in3 => \N__33932\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34094\,
            in2 => \_gnd_net_\,
            in3 => \N__34085\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34082\,
            in2 => \_gnd_net_\,
            in3 => \N__34073\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34109\,
            in2 => \_gnd_net_\,
            in3 => \N__34070\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34067\,
            in2 => \_gnd_net_\,
            in3 => \N__34058\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34055\,
            in2 => \_gnd_net_\,
            in3 => \N__34046\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34043\,
            in2 => \_gnd_net_\,
            in3 => \N__34025\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34022\,
            in2 => \_gnd_net_\,
            in3 => \N__34013\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34010\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39980\,
            in2 => \N__33995\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38793\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__38512\,
            in1 => \N__38489\,
            in2 => \_gnd_net_\,
            in3 => \N__40107\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40110\,
            in1 => \N__38549\,
            in2 => \_gnd_net_\,
            in3 => \N__38525\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38309\,
            in1 => \N__40109\,
            in2 => \_gnd_net_\,
            in3 => \N__38279\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38383\,
            in1 => \N__40108\,
            in2 => \_gnd_net_\,
            in3 => \N__38357\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38259\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38508\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34103\,
            ce => 'H',
            sr => \N__44182\
        );

    \delay_measurement_inst.start_timer_tr_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36714\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34103\,
            ce => 'H',
            sr => \N__44182\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__34478\,
            in1 => \N__34454\,
            in2 => \N__34962\,
            in3 => \N__34424\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34385\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34324\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34566\,
            in2 => \_gnd_net_\,
            in3 => \N__35079\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35149\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34631\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35306\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35737\,
            in1 => \N__35648\,
            in2 => \N__35512\,
            in3 => \N__34253\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44931\,
            ce => 'H',
            sr => \N__44109\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__35736\,
            in1 => \N__34247\,
            in2 => \_gnd_net_\,
            in3 => \N__34193\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__35646\,
            in1 => \N__35740\,
            in2 => \N__35515\,
            in3 => \N__35237\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44931\,
            ce => 'H',
            sr => \N__44109\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35738\,
            in1 => \N__35649\,
            in2 => \N__35513\,
            in3 => \N__35180\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44931\,
            ce => 'H',
            sr => \N__44109\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__35647\,
            in1 => \N__35741\,
            in2 => \N__35516\,
            in3 => \N__35120\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44931\,
            ce => 'H',
            sr => \N__44109\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35739\,
            in1 => \N__35650\,
            in2 => \N__35514\,
            in3 => \N__35063\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44931\,
            ce => 'H',
            sr => \N__44109\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__34630\,
            in1 => \N__34994\,
            in2 => \N__34963\,
            in3 => \N__34682\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__34658\,
            in1 => \N__35763\,
            in2 => \N__35673\,
            in3 => \N__35506\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44924\,
            ce => 'H',
            sr => \N__44114\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35759\,
            in1 => \N__35653\,
            in2 => \N__35518\,
            in3 => \N__34601\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44924\,
            ce => 'H',
            sr => \N__44114\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35651\,
            in1 => \N__35761\,
            in2 => \N__34544\,
            in3 => \N__35504\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44924\,
            ce => 'H',
            sr => \N__44114\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35760\,
            in1 => \N__35654\,
            in2 => \N__35519\,
            in3 => \N__35900\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44924\,
            ce => 'H',
            sr => \N__44114\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__35891\,
            in1 => \N__35762\,
            in2 => \N__35674\,
            in3 => \N__35505\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44924\,
            ce => 'H',
            sr => \N__44114\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__35758\,
            in1 => \N__35652\,
            in2 => \N__35517\,
            in3 => \N__35339\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44924\,
            ce => 'H',
            sr => \N__44114\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36009\,
            in1 => \N__38671\,
            in2 => \N__38650\,
            in3 => \N__35251\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__38646\,
            in1 => \N__39157\,
            in2 => \N__39184\,
            in3 => \N__36010\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__39234\,
            in1 => \N__35258\,
            in2 => \N__35276\,
            in3 => \N__35252\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38873\,
            in1 => \N__39204\,
            in2 => \N__39004\,
            in3 => \N__38571\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__38596\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38620\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39177\,
            in1 => \N__39156\,
            in2 => \N__39238\,
            in3 => \N__39205\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_367\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38572\,
            in1 => \N__38874\,
            in2 => \N__36044\,
            in3 => \N__38999\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__40750\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44918\,
            ce => \N__39291\,
            sr => \N__44118\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__39000\,
            in1 => \N__35933\,
            in2 => \_gnd_net_\,
            in3 => \N__35939\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__39452\,
            in1 => \N__35990\,
            in2 => \N__36547\,
            in3 => \N__36124\,
            lcout => \elapsed_time_ns_1_RNIVEIF91_0_25\,
            ltout => \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_o5_6_15_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35971\,
            in1 => \N__36193\,
            in2 => \N__35984\,
            in3 => \N__36232\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_i_o5_6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__36529\,
            in1 => \N__39410\,
            in2 => \N__35975\,
            in3 => \N__36125\,
            lcout => \elapsed_time_ns_1_RNI2IIF91_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__39060\,
            in1 => \N__38570\,
            in2 => \N__39037\,
            in3 => \N__35950\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38926\,
            in1 => \N__38947\,
            in2 => \N__38908\,
            in3 => \N__38968\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_347\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39061\,
            in1 => \N__39261\,
            in2 => \N__35927\,
            in3 => \N__39033\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36698\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39451\,
            in1 => \N__39130\,
            in2 => \N__39437\,
            in3 => \N__36221\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39361\,
            in1 => \N__39406\,
            in2 => \N__39388\,
            in3 => \N__39421\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__39436\,
            in1 => \N__36236\,
            in2 => \N__36554\,
            in3 => \N__36128\,
            lcout => \elapsed_time_ns_1_RNI0GIF91_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39112\,
            in1 => \N__39478\,
            in2 => \N__39091\,
            in3 => \N__39466\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__39479\,
            in1 => \N__36126\,
            in2 => \N__36215\,
            in3 => \N__36548\,
            lcout => \elapsed_time_ns_1_RNITCIF91_0_23\,
            ltout => \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_15_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36055\,
            in2 => \N__36206\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__36127\,
            in1 => \N__39422\,
            in2 => \N__36197\,
            in3 => \N__36549\,
            lcout => \elapsed_time_ns_1_RNI1HIF91_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__39467\,
            in1 => \N__36502\,
            in2 => \N__36059\,
            in3 => \N__36129\,
            lcout => \elapsed_time_ns_1_RNIUDIF91_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__36696\,
            in1 => \N__36724\,
            in2 => \_gnd_net_\,
            in3 => \N__36673\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_435_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__36674\,
            in1 => \_gnd_net_\,
            in2 => \N__36728\,
            in3 => \N__36697\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44906\,
            ce => 'H',
            sr => \N__44125\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36692\,
            in2 => \_gnd_net_\,
            in3 => \N__36672\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_434_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36631\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36596\,
            lcout => \phase_controller_inst1.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__41551\,
            in1 => \N__36525\,
            in2 => \N__38888\,
            in3 => \N__36377\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36329\,
            in3 => \N__36326\,
            lcout => \elapsed_time_ns_1_RNIDE4DM1_0_14\,
            ltout => \elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_6_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37018\,
            in2 => \N__36269\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_8_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__37586\,
            in1 => \N__42197\,
            in2 => \_gnd_net_\,
            in3 => \N__36837\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44901\,
            ce => \N__43745\,
            sr => \N__44129\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_7_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__42196\,
            in1 => \N__36871\,
            in2 => \_gnd_net_\,
            in3 => \N__37585\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44901\,
            ce => \N__43745\,
            sr => \N__44129\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a0_6_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__37019\,
            in1 => \N__36926\,
            in2 => \_gnd_net_\,
            in3 => \N__36899\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_0_6_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__36969\,
            in1 => \N__36887\,
            in2 => \N__36881\,
            in3 => \N__42025\,
            lcout => \phase_controller_inst1.stoper_tr.N_249\,
            ltout => \phase_controller_inst1.stoper_tr.N_249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_6_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__36813\,
            in1 => \N__42198\,
            in2 => \N__36878\,
            in3 => \N__36776\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44901\,
            ce => \N__43745\,
            sr => \N__44129\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_9_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__37195\,
            in1 => \N__42038\,
            in2 => \N__37217\,
            in3 => \N__42194\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44895\,
            ce => \N__41934\,
            sr => \N__44131\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_12_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__42187\,
            in1 => \N__42429\,
            in2 => \N__42074\,
            in3 => \N__41596\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44895\,
            ce => \N__41934\,
            sr => \N__44131\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_15_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__36970\,
            in1 => \N__42190\,
            in2 => \N__37033\,
            in3 => \N__42042\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44895\,
            ce => \N__41934\,
            sr => \N__44131\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_7_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__42186\,
            in1 => \_gnd_net_\,
            in2 => \N__36875\,
            in3 => \N__37588\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44895\,
            ce => \N__41934\,
            sr => \N__44131\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_8_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__37589\,
            in1 => \N__42189\,
            in2 => \_gnd_net_\,
            in3 => \N__36842\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44895\,
            ce => \N__41934\,
            sr => \N__44131\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_6_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__36814\,
            in1 => \N__37587\,
            in2 => \N__42227\,
            in3 => \N__36774\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44895\,
            ce => \N__41934\,
            sr => \N__44131\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_2_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001110"
        )
    port map (
            in0 => \N__37590\,
            in1 => \N__37488\,
            in2 => \N__37049\,
            in3 => \N__42195\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44895\,
            ce => \N__41934\,
            sr => \N__44131\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_5_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__42188\,
            in1 => \N__37591\,
            in2 => \N__37497\,
            in3 => \N__36943\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44895\,
            ce => \N__41934\,
            sr => \N__44131\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_9_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__42179\,
            in1 => \N__37216\,
            in2 => \N__37199\,
            in3 => \N__42073\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44890\,
            ce => \N__43735\,
            sr => \N__44139\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_17_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__42070\,
            in1 => \N__42304\,
            in2 => \_gnd_net_\,
            in3 => \N__42185\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44890\,
            ce => \N__43735\,
            sr => \N__44139\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_16_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__42180\,
            in1 => \N__42500\,
            in2 => \_gnd_net_\,
            in3 => \N__42072\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44890\,
            ce => \N__43735\,
            sr => \N__44139\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0_2_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010101"
        )
    port map (
            in0 => \N__37181\,
            in1 => \N__37153\,
            in2 => \N__37127\,
            in3 => \N__37087\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_2_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001100"
        )
    port map (
            in0 => \N__42181\,
            in1 => \N__37493\,
            in2 => \N__37040\,
            in3 => \N__37616\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44890\,
            ce => \N__43735\,
            sr => \N__44139\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_15_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__42071\,
            in1 => \N__42183\,
            in2 => \N__37037\,
            in3 => \N__36977\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44890\,
            ce => \N__43735\,
            sr => \N__44139\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_5_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__42182\,
            in1 => \N__36947\,
            in2 => \N__37498\,
            in3 => \N__37618\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44890\,
            ce => \N__43735\,
            sr => \N__44139\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_4_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__37617\,
            in1 => \N__42184\,
            in2 => \N__37544\,
            in3 => \N__37492\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44890\,
            ce => \N__43735\,
            sr => \N__44139\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__37698\,
            in1 => \N__37457\,
            in2 => \_gnd_net_\,
            in3 => \N__37435\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_c_RNO_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40003\,
            in1 => \N__37808\,
            in2 => \_gnd_net_\,
            in3 => \N__37778\,
            lcout => \current_shift_inst.un38_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__37695\,
            in1 => \N__37411\,
            in2 => \_gnd_net_\,
            in3 => \N__37399\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__37375\,
            in1 => \N__37699\,
            in2 => \_gnd_net_\,
            in3 => \N__37351\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__37701\,
            in1 => \N__37340\,
            in2 => \_gnd_net_\,
            in3 => \N__37312\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__37301\,
            in1 => \N__37696\,
            in2 => \_gnd_net_\,
            in3 => \N__37270\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__37697\,
            in1 => \N__37258\,
            in2 => \_gnd_net_\,
            in3 => \N__37228\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__37975\,
            in1 => \N__37700\,
            in2 => \_gnd_net_\,
            in3 => \N__37945\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__37933\,
            in1 => \N__37720\,
            in2 => \_gnd_net_\,
            in3 => \N__37903\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__37723\,
            in1 => \N__37892\,
            in2 => \_gnd_net_\,
            in3 => \N__37864\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37833\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__37725\,
            in1 => \N__38029\,
            in2 => \_gnd_net_\,
            in3 => \N__38002\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__37846\,
            in1 => \N__37726\,
            in2 => \_gnd_net_\,
            in3 => \N__37834\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__37722\,
            in1 => \N__37807\,
            in2 => \_gnd_net_\,
            in3 => \N__37777\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__37766\,
            in1 => \N__37724\,
            in2 => \_gnd_net_\,
            in3 => \N__37741\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__37721\,
            in1 => \N__37661\,
            in2 => \_gnd_net_\,
            in3 => \N__37633\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38156\,
            in1 => \N__39963\,
            in2 => \_gnd_net_\,
            in3 => \N__38132\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38203\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44870\,
            ce => \N__38179\,
            sr => \N__44157\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38155\,
            in1 => \N__39961\,
            in2 => \_gnd_net_\,
            in3 => \N__38131\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__39957\,
            in1 => \N__38074\,
            in2 => \_gnd_net_\,
            in3 => \N__38065\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__38747\,
            in1 => \N__38710\,
            in2 => \_gnd_net_\,
            in3 => \N__39958\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39959\,
            in1 => \N__38122\,
            in2 => \_gnd_net_\,
            in3 => \N__38086\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38800\,
            in1 => \N__39960\,
            in2 => \_gnd_net_\,
            in3 => \N__38770\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_c_RNO_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__39962\,
            in1 => \N__38075\,
            in2 => \_gnd_net_\,
            in3 => \N__38066\,
            lcout => \current_shift_inst.un38_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_c_RNO_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38033\,
            in1 => \N__39978\,
            in2 => \_gnd_net_\,
            in3 => \N__38006\,
            lcout => \current_shift_inst.un38_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39977\,
            in1 => \N__38548\,
            in2 => \_gnd_net_\,
            in3 => \N__38524\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38513\,
            in1 => \N__39974\,
            in2 => \_gnd_net_\,
            in3 => \N__38488\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_c_RNO_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39979\,
            in1 => \N__38477\,
            in2 => \_gnd_net_\,
            in3 => \N__38459\,
            lcout => \current_shift_inst.un38_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38431\,
            in1 => \N__39976\,
            in2 => \_gnd_net_\,
            in3 => \N__38395\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39973\,
            in1 => \N__38384\,
            in2 => \_gnd_net_\,
            in3 => \N__38353\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38342\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39975\,
            in1 => \N__38308\,
            in2 => \_gnd_net_\,
            in3 => \N__38278\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39995\,
            in1 => \N__38267\,
            in2 => \_gnd_net_\,
            in3 => \N__38237\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__39999\,
            in1 => \N__38819\,
            in2 => \_gnd_net_\,
            in3 => \N__38840\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38839\,
            in1 => \N__39996\,
            in2 => \_gnd_net_\,
            in3 => \N__38818\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38804\,
            in1 => \N__39998\,
            in2 => \_gnd_net_\,
            in3 => \N__38774\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_c_RNO_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__39997\,
            in1 => \N__38746\,
            in2 => \_gnd_net_\,
            in3 => \N__38717\,
            lcout => \current_shift_inst.un38_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40778\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44932\,
            ce => \N__39292\,
            sr => \N__44110\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40777\,
            in2 => \N__40720\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__44925\,
            ce => \N__39293\,
            sr => \N__44115\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40693\,
            in2 => \N__40751\,
            in3 => \N__38609\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__44925\,
            ce => \N__39293\,
            sr => \N__44115\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41065\,
            in2 => \N__40721\,
            in3 => \N__38585\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__44925\,
            ce => \N__39293\,
            sr => \N__44115\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40694\,
            in2 => \N__41036\,
            in3 => \N__38552\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__44925\,
            ce => \N__39293\,
            sr => \N__44115\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41005\,
            in2 => \N__41066\,
            in3 => \N__39047\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__44925\,
            ce => \N__39293\,
            sr => \N__44115\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41032\,
            in2 => \N__40984\,
            in3 => \N__39014\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__44925\,
            ce => \N__39293\,
            sr => \N__44115\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41006\,
            in2 => \N__40957\,
            in3 => \N__38978\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__44925\,
            ce => \N__39293\,
            sr => \N__44115\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40920\,
            in2 => \N__40985\,
            in3 => \N__38957\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__44925\,
            ce => \N__39293\,
            sr => \N__44115\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40958\,
            in2 => \N__40894\,
            in3 => \N__38936\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__44919\,
            ce => \N__39294\,
            sr => \N__44119\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40867\,
            in2 => \N__40928\,
            in3 => \N__38915\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__44919\,
            ce => \N__39294\,
            sr => \N__44119\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40846\,
            in2 => \N__40895\,
            in3 => \N__38891\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__44919\,
            ce => \N__39294\,
            sr => \N__44119\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40868\,
            in2 => \N__41285\,
            in3 => \N__38855\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__44919\,
            ce => \N__39294\,
            sr => \N__44119\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41254\,
            in2 => \N__40847\,
            in3 => \N__39248\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__44919\,
            ce => \N__39294\,
            sr => \N__44119\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41281\,
            in2 => \N__41233\,
            in3 => \N__39215\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__44919\,
            ce => \N__39294\,
            sr => \N__44119\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41255\,
            in2 => \N__41206\,
            in3 => \N__39191\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__44919\,
            ce => \N__39294\,
            sr => \N__44119\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41170\,
            in2 => \N__41234\,
            in3 => \N__39164\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__44919\,
            ce => \N__39294\,
            sr => \N__44119\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41207\,
            in2 => \N__41143\,
            in3 => \N__39137\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__44914\,
            ce => \N__39295\,
            sr => \N__44121\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41116\,
            in2 => \N__41177\,
            in3 => \N__39119\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__44914\,
            ce => \N__39295\,
            sr => \N__44121\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41095\,
            in2 => \N__41144\,
            in3 => \N__39095\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__44914\,
            ce => \N__39295\,
            sr => \N__44121\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41117\,
            in2 => \N__41495\,
            in3 => \N__39071\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__44914\,
            ce => \N__39295\,
            sr => \N__44121\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41464\,
            in2 => \N__41096\,
            in3 => \N__39470\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__44914\,
            ce => \N__39295\,
            sr => \N__44121\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41491\,
            in2 => \N__41443\,
            in3 => \N__39455\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__44914\,
            ce => \N__39295\,
            sr => \N__44121\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41465\,
            in2 => \N__41416\,
            in3 => \N__39440\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__44914\,
            ce => \N__39295\,
            sr => \N__44121\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41379\,
            in2 => \N__41444\,
            in3 => \N__39425\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__44914\,
            ce => \N__39295\,
            sr => \N__44121\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41417\,
            in2 => \N__41353\,
            in3 => \N__39413\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__44910\,
            ce => \N__39296\,
            sr => \N__44123\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41326\,
            in2 => \N__41387\,
            in3 => \N__39395\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__44910\,
            ce => \N__39296\,
            sr => \N__44123\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41306\,
            in2 => \N__41354\,
            in3 => \N__39371\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__44910\,
            ce => \N__39296\,
            sr => \N__44123\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41327\,
            in2 => \N__41678\,
            in3 => \N__39350\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__44910\,
            ce => \N__39296\,
            sr => \N__44123\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39347\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44910\,
            ce => \N__39296\,
            sr => \N__44123\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41888\,
            in2 => \N__39518\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41849\,
            in2 => \_gnd_net_\,
            in3 => \N__39503\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \N__44907\,
            ce => 'H',
            sr => \N__39664\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43106\,
            in2 => \N__42764\,
            in3 => \N__39500\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \N__44907\,
            ce => 'H',
            sr => \N__39664\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42728\,
            in2 => \_gnd_net_\,
            in3 => \N__39497\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \N__44907\,
            ce => 'H',
            sr => \N__39664\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42695\,
            in2 => \_gnd_net_\,
            in3 => \N__39494\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \N__44907\,
            ce => 'H',
            sr => \N__39664\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42662\,
            in2 => \_gnd_net_\,
            in3 => \N__39491\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \N__44907\,
            ce => 'H',
            sr => \N__39664\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42629\,
            in2 => \_gnd_net_\,
            in3 => \N__39488\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \N__44907\,
            ce => 'H',
            sr => \N__39664\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42605\,
            in2 => \_gnd_net_\,
            in3 => \N__39485\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \N__44907\,
            ce => 'H',
            sr => \N__39664\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42560\,
            in2 => \_gnd_net_\,
            in3 => \N__39482\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \N__44902\,
            ce => 'H',
            sr => \N__39657\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43031\,
            in2 => \_gnd_net_\,
            in3 => \N__39545\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \N__44902\,
            ce => 'H',
            sr => \N__39657\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42992\,
            in2 => \_gnd_net_\,
            in3 => \N__39542\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \N__44902\,
            ce => 'H',
            sr => \N__39657\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42959\,
            in2 => \_gnd_net_\,
            in3 => \N__39539\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \N__44902\,
            ce => 'H',
            sr => \N__39657\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42926\,
            in2 => \_gnd_net_\,
            in3 => \N__39536\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \N__44902\,
            ce => 'H',
            sr => \N__39657\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42896\,
            in2 => \_gnd_net_\,
            in3 => \N__39533\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \N__44902\,
            ce => 'H',
            sr => \N__39657\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42860\,
            in2 => \_gnd_net_\,
            in3 => \N__39530\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \N__44902\,
            ce => 'H',
            sr => \N__39657\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42842\,
            in2 => \_gnd_net_\,
            in3 => \N__39527\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \N__44902\,
            ce => 'H',
            sr => \N__39657\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42800\,
            in2 => \_gnd_net_\,
            in3 => \N__39524\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \N__44896\,
            ce => 'H',
            sr => \N__39665\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43253\,
            in2 => \_gnd_net_\,
            in3 => \N__39521\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \N__44896\,
            ce => 'H',
            sr => \N__39665\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43214\,
            in2 => \_gnd_net_\,
            in3 => \N__39668\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44896\,
            ce => 'H',
            sr => \N__39665\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39623\,
            in2 => \N__39611\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40594\,
            in2 => \N__39596\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39581\,
            in2 => \N__40620\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40598\,
            in2 => \N__39575\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39566\,
            in2 => \N__40621\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40602\,
            in2 => \N__39560\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39551\,
            in2 => \N__40622\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40606\,
            in2 => \N__39740\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40590\,
            in2 => \N__39728\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39719\,
            in2 => \N__40619\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40578\,
            in2 => \N__39713\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39704\,
            in2 => \N__40616\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40582\,
            in2 => \N__39698\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39689\,
            in2 => \N__40617\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40586\,
            in2 => \N__39683\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39674\,
            in2 => \N__40618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39809\,
            in2 => \N__40574\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40502\,
            in2 => \N__39800\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39791\,
            in2 => \N__40575\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40506\,
            in2 => \N__39785\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39776\,
            in2 => \N__40576\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40510\,
            in2 => \N__39770\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39761\,
            in2 => \N__40577\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40514\,
            in2 => \N__39752\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40486\,
            in2 => \N__40673\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40664\,
            in2 => \N__40571\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40490\,
            in2 => \N__40658\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40649\,
            in2 => \N__40572\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40494\,
            in2 => \N__40643\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40628\,
            in2 => \N__40573\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40498\,
            in2 => \N__40292\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39991\,
            in2 => \_gnd_net_\,
            in3 => \N__39869\,
            lcout => \current_shift_inst.N_1310_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_RNIOA7T_1_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101110"
        )
    port map (
            in0 => \N__44320\,
            in1 => \N__43778\,
            in2 => \N__43832\,
            in3 => \N__43856\,
            lcout => \phase_controller_inst2.stoper_tr.un1_stoper_state12_1_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_0_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__43779\,
            in1 => \N__43819\,
            in2 => \N__43864\,
            in3 => \N__44380\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44864\,
            ce => 'H',
            sr => \N__44161\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43855\,
            in2 => \_gnd_net_\,
            in3 => \N__43777\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_tr.N_45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011001010"
        )
    port map (
            in0 => \N__43826\,
            in1 => \N__40800\,
            in2 => \N__40817\,
            in3 => \N__44381\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44864\,
            ce => 'H',
            sr => \N__44161\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_1_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__44379\,
            in1 => \N__43780\,
            in2 => \N__43833\,
            in3 => \N__43860\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44864\,
            ce => 'H',
            sr => \N__44161\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41814\,
            in1 => \N__40765\,
            in2 => \_gnd_net_\,
            in3 => \N__40754\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__44941\,
            ce => \N__41657\,
            sr => \N__44103\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41809\,
            in1 => \N__40740\,
            in2 => \_gnd_net_\,
            in3 => \N__40724\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__44941\,
            ce => \N__41657\,
            sr => \N__44103\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41815\,
            in1 => \N__40713\,
            in2 => \_gnd_net_\,
            in3 => \N__40697\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__44941\,
            ce => \N__41657\,
            sr => \N__44103\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41810\,
            in1 => \N__40692\,
            in2 => \_gnd_net_\,
            in3 => \N__40676\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__44941\,
            ce => \N__41657\,
            sr => \N__44103\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41816\,
            in1 => \N__41058\,
            in2 => \_gnd_net_\,
            in3 => \N__41039\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__44941\,
            ce => \N__41657\,
            sr => \N__44103\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41811\,
            in1 => \N__41028\,
            in2 => \_gnd_net_\,
            in3 => \N__41009\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__44941\,
            ce => \N__41657\,
            sr => \N__44103\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41813\,
            in1 => \N__41004\,
            in2 => \_gnd_net_\,
            in3 => \N__40988\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__44941\,
            ce => \N__41657\,
            sr => \N__44103\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41812\,
            in1 => \N__40977\,
            in2 => \_gnd_net_\,
            in3 => \N__40961\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__44941\,
            ce => \N__41657\,
            sr => \N__44103\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41798\,
            in1 => \N__40950\,
            in2 => \_gnd_net_\,
            in3 => \N__40931\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__44938\,
            ce => \N__41656\,
            sr => \N__44104\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41794\,
            in1 => \N__40924\,
            in2 => \_gnd_net_\,
            in3 => \N__40898\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__44938\,
            ce => \N__41656\,
            sr => \N__44104\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41795\,
            in1 => \N__40887\,
            in2 => \_gnd_net_\,
            in3 => \N__40871\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__44938\,
            ce => \N__41656\,
            sr => \N__44104\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41791\,
            in1 => \N__40866\,
            in2 => \_gnd_net_\,
            in3 => \N__40850\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__44938\,
            ce => \N__41656\,
            sr => \N__44104\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41796\,
            in1 => \N__40839\,
            in2 => \_gnd_net_\,
            in3 => \N__40820\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__44938\,
            ce => \N__41656\,
            sr => \N__44104\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41792\,
            in1 => \N__41277\,
            in2 => \_gnd_net_\,
            in3 => \N__41258\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__44938\,
            ce => \N__41656\,
            sr => \N__44104\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41797\,
            in1 => \N__41253\,
            in2 => \_gnd_net_\,
            in3 => \N__41237\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__44938\,
            ce => \N__41656\,
            sr => \N__44104\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41793\,
            in1 => \N__41226\,
            in2 => \_gnd_net_\,
            in3 => \N__41210\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__44938\,
            ce => \N__41656\,
            sr => \N__44104\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41787\,
            in1 => \N__41199\,
            in2 => \_gnd_net_\,
            in3 => \N__41180\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_18_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__44935\,
            ce => \N__41655\,
            sr => \N__44106\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41803\,
            in1 => \N__41169\,
            in2 => \_gnd_net_\,
            in3 => \N__41147\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__44935\,
            ce => \N__41655\,
            sr => \N__44106\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41788\,
            in1 => \N__41136\,
            in2 => \_gnd_net_\,
            in3 => \N__41120\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__44935\,
            ce => \N__41655\,
            sr => \N__44106\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41804\,
            in1 => \N__41115\,
            in2 => \_gnd_net_\,
            in3 => \N__41099\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__44935\,
            ce => \N__41655\,
            sr => \N__44106\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41789\,
            in1 => \N__41088\,
            in2 => \_gnd_net_\,
            in3 => \N__41069\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__44935\,
            ce => \N__41655\,
            sr => \N__44106\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41805\,
            in1 => \N__41487\,
            in2 => \_gnd_net_\,
            in3 => \N__41468\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__44935\,
            ce => \N__41655\,
            sr => \N__44106\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41790\,
            in1 => \N__41463\,
            in2 => \_gnd_net_\,
            in3 => \N__41447\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__44935\,
            ce => \N__41655\,
            sr => \N__44106\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41806\,
            in1 => \N__41436\,
            in2 => \_gnd_net_\,
            in3 => \N__41420\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__44935\,
            ce => \N__41655\,
            sr => \N__44106\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41799\,
            in1 => \N__41409\,
            in2 => \_gnd_net_\,
            in3 => \N__41390\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__44933\,
            ce => \N__41645\,
            sr => \N__44111\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41807\,
            in1 => \N__41383\,
            in2 => \_gnd_net_\,
            in3 => \N__41357\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__44933\,
            ce => \N__41645\,
            sr => \N__44111\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41800\,
            in1 => \N__41346\,
            in2 => \_gnd_net_\,
            in3 => \N__41330\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__44933\,
            ce => \N__41645\,
            sr => \N__44111\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41808\,
            in1 => \N__41325\,
            in2 => \_gnd_net_\,
            in3 => \N__41309\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__44933\,
            ce => \N__41645\,
            sr => \N__44111\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41801\,
            in1 => \N__41302\,
            in2 => \_gnd_net_\,
            in3 => \N__41288\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__44933\,
            ce => \N__41645\,
            sr => \N__44111\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__41671\,
            in1 => \N__41802\,
            in2 => \_gnd_net_\,
            in3 => \N__41681\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44933\,
            ce => \N__41645\,
            sr => \N__44111\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_14_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__41567\,
            in1 => \N__42266\,
            in2 => \N__42089\,
            in3 => \N__42454\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44926\,
            ce => \N__43744\,
            sr => \N__44116\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_10_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__42450\,
            in1 => \N__42067\,
            in2 => \N__42269\,
            in3 => \N__41527\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44926\,
            ce => \N__43744\,
            sr => \N__44116\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_11_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__42061\,
            in1 => \N__42264\,
            in2 => \N__42539\,
            in3 => \N__42452\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44926\,
            ce => \N__43744\,
            sr => \N__44116\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_13_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__42062\,
            in1 => \N__42265\,
            in2 => \N__42413\,
            in3 => \N__42453\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44926\,
            ce => \N__43744\,
            sr => \N__44116\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_12_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__42451\,
            in1 => \N__42256\,
            in2 => \N__41600\,
            in3 => \N__42068\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44926\,
            ce => \N__43744\,
            sr => \N__44116\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_19_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__42060\,
            in1 => \_gnd_net_\,
            in2 => \N__42268\,
            in3 => \N__42380\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44926\,
            ce => \N__43744\,
            sr => \N__44116\
        );

    \phase_controller_inst2.stoper_tr.target_time_esr_18_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__42260\,
            in1 => \N__42343\,
            in2 => \_gnd_net_\,
            in3 => \N__42066\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44926\,
            ce => \N__43744\,
            sr => \N__44116\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_14_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__42457\,
            in1 => \N__41566\,
            in2 => \N__42092\,
            in3 => \N__42248\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44920\,
            ce => \N__41945\,
            sr => \N__44120\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_10_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__42244\,
            in1 => \N__42458\,
            in2 => \N__41528\,
            in3 => \N__42088\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44920\,
            ce => \N__41945\,
            sr => \N__44120\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_11_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__42455\,
            in1 => \N__42245\,
            in2 => \N__42090\,
            in3 => \N__42534\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44920\,
            ce => \N__41945\,
            sr => \N__44120\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_16_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__42494\,
            in1 => \N__42249\,
            in2 => \_gnd_net_\,
            in3 => \N__42085\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44920\,
            ce => \N__41945\,
            sr => \N__44120\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_13_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__42456\,
            in1 => \N__42246\,
            in2 => \N__42091\,
            in3 => \N__42412\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44920\,
            ce => \N__41945\,
            sr => \N__44120\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_19_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__42379\,
            in1 => \N__42251\,
            in2 => \_gnd_net_\,
            in3 => \N__42087\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44920\,
            ce => \N__41945\,
            sr => \N__44120\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_18_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__42075\,
            in1 => \N__42344\,
            in2 => \_gnd_net_\,
            in3 => \N__42247\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44920\,
            ce => \N__41945\,
            sr => \N__44120\
        );

    \phase_controller_inst1.stoper_tr.target_time_esr_17_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__42305\,
            in1 => \N__42250\,
            in2 => \_gnd_net_\,
            in3 => \N__42086\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44920\,
            ce => \N__41945\,
            sr => \N__44120\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41906\,
            in2 => \N__41861\,
            in3 => \N__41881\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__41848\,
            in1 => \N__41837\,
            in2 => \N__41825\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42749\,
            in2 => \N__42782\,
            in3 => \N__42760\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42743\,
            in2 => \N__42716\,
            in3 => \N__42727\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42707\,
            in2 => \N__42683\,
            in3 => \N__42694\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42674\,
            in2 => \N__42650\,
            in3 => \N__42661\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42641\,
            in2 => \N__42617\,
            in3 => \N__42628\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__42604\,
            in1 => \N__42593\,
            in2 => \N__42581\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42572\,
            in2 => \N__42548\,
            in3 => \N__42559\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43030\,
            in1 => \N__43019\,
            in2 => \N__43010\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43001\,
            in2 => \N__42980\,
            in3 => \N__42991\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42971\,
            in2 => \N__42947\,
            in3 => \N__42958\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42914\,
            in2 => \N__42938\,
            in3 => \N__42925\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42905\,
            in2 => \N__42884\,
            in3 => \N__42895\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42848\,
            in2 => \N__42875\,
            in3 => \N__42859\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__42841\,
            in1 => \N__42830\,
            in2 => \N__42821\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42788\,
            in2 => \N__42812\,
            in3 => \N__42799\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43252\,
            in1 => \N__43241\,
            in2 => \N__43232\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43223\,
            in2 => \N__43202\,
            in3 => \N__43213\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43193\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NA_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43189\,
            in2 => \_gnd_net_\,
            in3 => \N__43131\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43085\,
            in2 => \N__43100\,
            in3 => \N__43681\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43079\,
            in2 => \N__43070\,
            in3 => \N__43637\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43061\,
            in2 => \N__43049\,
            in3 => \N__43607\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43040\,
            in2 => \N__43406\,
            in3 => \N__43589\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43385\,
            in2 => \N__43397\,
            in3 => \N__44546\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44528\,
            in1 => \N__43379\,
            in2 => \N__43367\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43358\,
            in2 => \N__43346\,
            in3 => \N__44510\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43337\,
            in2 => \N__43325\,
            in3 => \N__44492\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43313\,
            in2 => \N__43298\,
            in3 => \N__44474\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43289\,
            in2 => \N__43280\,
            in3 => \N__44456\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43259\,
            in2 => \N__43271\,
            in3 => \N__44438\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43571\,
            in2 => \N__43559\,
            in3 => \N__44420\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43550\,
            in2 => \N__43538\,
            in3 => \N__44402\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45059\,
            in1 => \N__43529\,
            in2 => \N__43520\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43511\,
            in2 => \N__43499\,
            in3 => \N__45041\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43475\,
            in2 => \N__43490\,
            in3 => \N__45023\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43469\,
            in2 => \N__43457\,
            in3 => \N__45005\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43448\,
            in2 => \N__43439\,
            in3 => \N__44987\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43427\,
            in2 => \N__43415\,
            in3 => \N__44966\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44384\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84AD_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__43828\,
            in1 => \_gnd_net_\,
            in2 => \N__44367\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84ADZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43827\,
            in2 => \_gnd_net_\,
            in3 => \N__44357\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_RNIOA7T_0_1_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__44315\,
            in1 => \N__43868\,
            in2 => \N__43837\,
            in3 => \N__43784\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43682\,
            in2 => \N__43646\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43636\,
            in2 => \_gnd_net_\,
            in3 => \N__43622\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \N__44885\,
            ce => 'H',
            sr => \N__44587\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43606\,
            in2 => \N__43619\,
            in3 => \N__43592\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \N__44885\,
            ce => 'H',
            sr => \N__44587\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43588\,
            in2 => \_gnd_net_\,
            in3 => \N__43574\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \N__44885\,
            ce => 'H',
            sr => \N__44587\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44545\,
            in2 => \_gnd_net_\,
            in3 => \N__44531\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \N__44885\,
            ce => 'H',
            sr => \N__44587\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44527\,
            in2 => \_gnd_net_\,
            in3 => \N__44513\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \N__44885\,
            ce => 'H',
            sr => \N__44587\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44509\,
            in2 => \_gnd_net_\,
            in3 => \N__44495\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \N__44885\,
            ce => 'H',
            sr => \N__44587\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44491\,
            in2 => \_gnd_net_\,
            in3 => \N__44477\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \N__44885\,
            ce => 'H',
            sr => \N__44587\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44473\,
            in2 => \_gnd_net_\,
            in3 => \N__44459\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \N__44877\,
            ce => 'H',
            sr => \N__44577\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44455\,
            in2 => \_gnd_net_\,
            in3 => \N__44441\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \N__44877\,
            ce => 'H',
            sr => \N__44577\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44437\,
            in2 => \_gnd_net_\,
            in3 => \N__44423\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \N__44877\,
            ce => 'H',
            sr => \N__44577\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44419\,
            in2 => \_gnd_net_\,
            in3 => \N__44405\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \N__44877\,
            ce => 'H',
            sr => \N__44577\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44401\,
            in2 => \_gnd_net_\,
            in3 => \N__44387\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \N__44877\,
            ce => 'H',
            sr => \N__44577\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45058\,
            in2 => \_gnd_net_\,
            in3 => \N__45044\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \N__44877\,
            ce => 'H',
            sr => \N__44577\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45040\,
            in2 => \_gnd_net_\,
            in3 => \N__45026\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \N__44877\,
            ce => 'H',
            sr => \N__44577\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45022\,
            in2 => \_gnd_net_\,
            in3 => \N__45008\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \N__44877\,
            ce => 'H',
            sr => \N__44577\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45004\,
            in2 => \_gnd_net_\,
            in3 => \N__44990\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_18_21_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \N__44871\,
            ce => 'H',
            sr => \N__44576\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44986\,
            in2 => \_gnd_net_\,
            in3 => \N__44972\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \N__44871\,
            ce => 'H',
            sr => \N__44576\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44965\,
            in2 => \_gnd_net_\,
            in3 => \N__44969\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__44871\,
            ce => 'H',
            sr => \N__44576\
        );
end \INTERFACE\;
