-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 24 2025 22:19:58

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T45 : out std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    T01 : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__47639\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47592\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47529\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47500\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47491\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47338\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47177\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47104\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46948\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46618\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46130\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46103\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45601\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45109\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44993\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44747\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44290\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43782\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43307\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43049\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42541\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42410\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42386\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42292\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41906\ : std_logic;
signal \N__41903\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \rgb_drv_RNOZ0\ : std_logic;
signal \N_38_i_i\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \bfn_3_8_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_153\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_154\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \N_19_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\ : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_155\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_149\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_53\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74_16_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_72\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_1_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_432_i\ : std_logic;
signal il_max_comp1_c : std_logic;
signal il_max_comp2_c : std_logic;
signal il_min_comp2_c : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_62\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI3VBED1_0_16_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNI40CED1_0_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal il_min_comp1_c : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_275_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_325_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIB4DJ11_0_5_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIL13KD1_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_266_iZ0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNI3VBED1_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_287\ : std_logic;
signal \elapsed_time_ns_1_RNI1TBED1_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI51CED1_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI40CED1_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI62CED1_0_19\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal s3_phy_c : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_30\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIP1MD11_0_12_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_337\ : std_logic;
signal \elapsed_time_ns_1_RNINVLD11_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIP2ND11_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNIP2ND11_0_21_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIU7ND11_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNIR4ND11_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNIR4ND11_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNI0AND11_0_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNI1BND11_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNIO1ND11_0_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIV8ND11_0_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_10_25_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_10_26_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_103\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \elapsed_time_ns_1_RNIO0MD11_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIP1MD11_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10\ : std_logic;
signal \elapsed_time_ns_1_RNIQ2MD11_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNID6DJ11_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNIE7DJ11_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIDP2KD1_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_307\ : std_logic;
signal \elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNIA3DJ11_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_325\ : std_logic;
signal \elapsed_time_ns_1_RNIQ4OD11_0_31\ : std_logic;
signal \elapsed_time_ns_1_RNIB4DJ11_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_327\ : std_logic;
signal \elapsed_time_ns_1_RNIP3OD11_0_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_382_i_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIS5ND11_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNIT6ND11_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNIS4MD11_0_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNIQ3ND11_0_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIQURR91_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNIQURR91_0_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_283\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal s4_phy_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.N_55\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \phase_controller_inst1.N_56\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3DZ0Z41\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\ : std_logic;
signal \elapsed_time_ns_1_RNIIU2KD1_0_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5\ : std_logic;
signal \elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_12_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.time_passed_RNI9M3O_cascade_\ : std_logic;
signal state_3 : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_433_i\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.N_166_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIUKL2M1_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\ : std_logic;
signal \elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_211_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNIPFL2M1_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNICG2591_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNICG2591_0_4_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIFG4DM1_0_16\ : std_logic;
signal \elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIGH4DM1_0_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_251\ : std_logic;
signal \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNI1OL2M1_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6NZ0Z32\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_0_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_432_i_g\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_434_i\ : std_logic;
signal \bfn_15_5_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_15_6_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \elapsed_time_ns_1_RNIGK2591_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIHI4DM1_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_214\ : std_logic;
signal \elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIUCHF91_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_241_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_RNOZ0Z_0\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_435_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\ : std_logic;
signal \elapsed_time_ns_1_RNIAE2591_0_2\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \T45_c\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.control_input_1_axb_0\ : std_logic;
signal \current_shift_inst.N_1572_i\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_0\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_1_cry_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_8\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_16_25_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_167_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_434_i_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_341\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIRHL2M1_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_381_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_358_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_381\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_348_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \elapsed_time_ns_1_RNIFJ2591_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNITCIF91_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIRAIF91_0_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \elapsed_time_ns_1_RNIDH2591_0_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_347\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \elapsed_time_ns_1_RNIQ8HF91_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIQ8HF91_0_11_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIR9HF91_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_244\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \elapsed_time_ns_1_RNI3JIF91_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI3JIF91_0_29_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNIDE4DM1_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \elapsed_time_ns_1_RNISAHF91_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_241\ : std_logic;
signal \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_13\ : std_logic;
signal \elapsed_time_ns_1_RNIIJ4DM1_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNISCJF91_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_19\ : std_logic;
signal start_stop_c : std_logic;
signal state_ns_i_a3_1 : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.N_166_i_g\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_382_i\ : std_logic;
signal \elapsed_time_ns_1_RNI81DJ11_0_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \T01_c\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \T12_c\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_367\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_349\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_363_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_380\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_365\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_345\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_359_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \elapsed_time_ns_1_RNIUDIF91_0_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \elapsed_time_ns_1_RNIVEIF91_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI0GIF91_0_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \elapsed_time_ns_1_RNI2IIF91_0_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_378\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIP7HF91_0_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \elapsed_time_ns_1_RNI1HIF91_0_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \elapsed_time_ns_1_RNISBIF91_0_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \elapsed_time_ns_1_RNIQ9IF91_0_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNIRBJF91_0_30\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.time_passed_RNI9M3O\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLHZ0Z1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un4_control_input_0_31\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \T23_c\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal \T01_wire\ : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal \T12_wire\ : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal \T45_wire\ : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    T01 <= \T01_wire\;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    T12 <= \T12_wire\;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    T45 <= \T45_wire\;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__20002\&\N__19995\&\N__20000\&\N__19994\&\N__20001\&\N__19993\&\N__20003\&\N__19990\&\N__19996\&\N__19989\&\N__19997\&\N__19991\&\N__19998\&\N__19992\&\N__19999\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__37809\&\N__37806\&'0'&'0'&'0'&\N__37804\&\N__37808\&\N__37805\&\N__37807\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__20066\&\N__20045\&\N__20067\&\N__20046\&\N__20068\&\N__20456\&\N__20378\&\N__20416\&\N__20405\&\N__20284\&\N__20328\&\N__20354\&\N__19913\&\N__19886\&\N__19658\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__37729\&\N__37726\&'0'&'0'&'0'&\N__37724\&\N__37728\&\N__37725\&\N__37727\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__21362\,
            RESETB => \N__31034\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__37810\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__37803\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__37730\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__37723\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__47637\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47639\,
            DIN => \N__47638\,
            DOUT => \N__47637\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47639\,
            PADOUT => \N__47638\,
            PADIN => \N__47637\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T01_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47628\,
            DIN => \N__47627\,
            DOUT => \N__47626\,
            PACKAGEPIN => \T01_wire\
        );

    \T01_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47628\,
            PADOUT => \N__47627\,
            PADIN => \N__47626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__41909\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47619\,
            DIN => \N__47618\,
            DOUT => \N__47617\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47619\,
            PADOUT => \N__47618\,
            PADIN => \N__47617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47610\,
            DIN => \N__47609\,
            DOUT => \N__47608\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47610\,
            PADOUT => \N__47609\,
            PADIN => \N__47608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47601\,
            DIN => \N__47600\,
            DOUT => \N__47599\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47601\,
            PADOUT => \N__47600\,
            PADIN => \N__47599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__46133\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47592\,
            DIN => \N__47591\,
            DOUT => \N__47590\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47592\,
            PADOUT => \N__47591\,
            PADIN => \N__47590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22349\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47583\,
            DIN => \N__47582\,
            DOUT => \N__47581\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47583\,
            PADOUT => \N__47582\,
            PADIN => \N__47581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47574\,
            DIN => \N__47573\,
            DOUT => \N__47572\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47574\,
            PADOUT => \N__47573\,
            PADIN => \N__47572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31046\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47565\,
            DIN => \N__47564\,
            DOUT => \N__47563\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47565\,
            PADOUT => \N__47564\,
            PADIN => \N__47563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__41804\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47556\,
            DIN => \N__47555\,
            DOUT => \N__47554\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47556\,
            PADOUT => \N__47555\,
            PADIN => \N__47554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47547\,
            DIN => \N__47546\,
            DOUT => \N__47545\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47547\,
            PADOUT => \N__47546\,
            PADIN => \N__47545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31211\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47538\,
            DIN => \N__47537\,
            DOUT => \N__47536\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47538\,
            PADOUT => \N__47537\,
            PADIN => \N__47536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28664\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47529\,
            DIN => \N__47528\,
            DOUT => \N__47527\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47529\,
            PADOUT => \N__47528\,
            PADIN => \N__47527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47520\,
            DIN => \N__47519\,
            DOUT => \N__47518\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47520\,
            PADOUT => \N__47519\,
            PADIN => \N__47518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23615\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T45_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47511\,
            DIN => \N__47510\,
            DOUT => \N__47509\,
            PACKAGEPIN => \T45_wire\
        );

    \T45_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47511\,
            PADOUT => \N__47510\,
            PADIN => \N__47509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36809\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47502\,
            DIN => \N__47501\,
            DOUT => \N__47500\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47502\,
            PADOUT => \N__47501\,
            PADIN => \N__47500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47493\,
            DIN => \N__47492\,
            DOUT => \N__47491\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47493\,
            PADOUT => \N__47492\,
            PADIN => \N__47491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11239\ : CascadeMux
    port map (
            O => \N__47474\,
            I => \N__47471\
        );

    \I__11238\ : InMux
    port map (
            O => \N__47471\,
            I => \N__47467\
        );

    \I__11237\ : InMux
    port map (
            O => \N__47470\,
            I => \N__47463\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__47467\,
            I => \N__47460\
        );

    \I__11235\ : InMux
    port map (
            O => \N__47466\,
            I => \N__47457\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__47463\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__11233\ : Odrv12
    port map (
            O => \N__47460\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__47457\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__11231\ : CascadeMux
    port map (
            O => \N__47450\,
            I => \N__47446\
        );

    \I__11230\ : InMux
    port map (
            O => \N__47449\,
            I => \N__47443\
        );

    \I__11229\ : InMux
    port map (
            O => \N__47446\,
            I => \N__47440\
        );

    \I__11228\ : LocalMux
    port map (
            O => \N__47443\,
            I => \N__47436\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__47440\,
            I => \N__47433\
        );

    \I__11226\ : InMux
    port map (
            O => \N__47439\,
            I => \N__47430\
        );

    \I__11225\ : Span4Mux_h
    port map (
            O => \N__47436\,
            I => \N__47424\
        );

    \I__11224\ : Span4Mux_h
    port map (
            O => \N__47433\,
            I => \N__47424\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__47430\,
            I => \N__47421\
        );

    \I__11222\ : InMux
    port map (
            O => \N__47429\,
            I => \N__47418\
        );

    \I__11221\ : Odrv4
    port map (
            O => \N__47424\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11220\ : Odrv4
    port map (
            O => \N__47421\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__47418\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11218\ : InMux
    port map (
            O => \N__47411\,
            I => \N__47408\
        );

    \I__11217\ : LocalMux
    port map (
            O => \N__47408\,
            I => \N__47405\
        );

    \I__11216\ : Span4Mux_h
    port map (
            O => \N__47405\,
            I => \N__47402\
        );

    \I__11215\ : Odrv4
    port map (
            O => \N__47402\,
            I => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\
        );

    \I__11214\ : InMux
    port map (
            O => \N__47399\,
            I => \N__47396\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__47396\,
            I => \N__47393\
        );

    \I__11212\ : Span4Mux_v
    port map (
            O => \N__47393\,
            I => \N__47390\
        );

    \I__11211\ : Odrv4
    port map (
            O => \N__47390\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__11210\ : InMux
    port map (
            O => \N__47387\,
            I => \N__47384\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__47384\,
            I => \N__47381\
        );

    \I__11208\ : Span4Mux_h
    port map (
            O => \N__47381\,
            I => \N__47378\
        );

    \I__11207\ : Span4Mux_h
    port map (
            O => \N__47378\,
            I => \N__47375\
        );

    \I__11206\ : Span4Mux_h
    port map (
            O => \N__47375\,
            I => \N__47372\
        );

    \I__11205\ : Odrv4
    port map (
            O => \N__47372\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__11204\ : InMux
    port map (
            O => \N__47369\,
            I => \N__47347\
        );

    \I__11203\ : InMux
    port map (
            O => \N__47368\,
            I => \N__47329\
        );

    \I__11202\ : InMux
    port map (
            O => \N__47367\,
            I => \N__47322\
        );

    \I__11201\ : InMux
    port map (
            O => \N__47366\,
            I => \N__47311\
        );

    \I__11200\ : InMux
    port map (
            O => \N__47365\,
            I => \N__47311\
        );

    \I__11199\ : InMux
    port map (
            O => \N__47364\,
            I => \N__47311\
        );

    \I__11198\ : InMux
    port map (
            O => \N__47363\,
            I => \N__47311\
        );

    \I__11197\ : InMux
    port map (
            O => \N__47362\,
            I => \N__47311\
        );

    \I__11196\ : InMux
    port map (
            O => \N__47361\,
            I => \N__47308\
        );

    \I__11195\ : InMux
    port map (
            O => \N__47360\,
            I => \N__47299\
        );

    \I__11194\ : InMux
    port map (
            O => \N__47359\,
            I => \N__47299\
        );

    \I__11193\ : InMux
    port map (
            O => \N__47358\,
            I => \N__47299\
        );

    \I__11192\ : InMux
    port map (
            O => \N__47357\,
            I => \N__47299\
        );

    \I__11191\ : InMux
    port map (
            O => \N__47356\,
            I => \N__47292\
        );

    \I__11190\ : InMux
    port map (
            O => \N__47355\,
            I => \N__47292\
        );

    \I__11189\ : InMux
    port map (
            O => \N__47354\,
            I => \N__47292\
        );

    \I__11188\ : InMux
    port map (
            O => \N__47353\,
            I => \N__47289\
        );

    \I__11187\ : InMux
    port map (
            O => \N__47352\,
            I => \N__47286\
        );

    \I__11186\ : InMux
    port map (
            O => \N__47351\,
            I => \N__47281\
        );

    \I__11185\ : InMux
    port map (
            O => \N__47350\,
            I => \N__47281\
        );

    \I__11184\ : LocalMux
    port map (
            O => \N__47347\,
            I => \N__47278\
        );

    \I__11183\ : InMux
    port map (
            O => \N__47346\,
            I => \N__47265\
        );

    \I__11182\ : InMux
    port map (
            O => \N__47345\,
            I => \N__47265\
        );

    \I__11181\ : InMux
    port map (
            O => \N__47344\,
            I => \N__47265\
        );

    \I__11180\ : InMux
    port map (
            O => \N__47343\,
            I => \N__47265\
        );

    \I__11179\ : InMux
    port map (
            O => \N__47342\,
            I => \N__47265\
        );

    \I__11178\ : InMux
    port map (
            O => \N__47341\,
            I => \N__47265\
        );

    \I__11177\ : InMux
    port map (
            O => \N__47340\,
            I => \N__47258\
        );

    \I__11176\ : InMux
    port map (
            O => \N__47339\,
            I => \N__47258\
        );

    \I__11175\ : InMux
    port map (
            O => \N__47338\,
            I => \N__47258\
        );

    \I__11174\ : InMux
    port map (
            O => \N__47337\,
            I => \N__47253\
        );

    \I__11173\ : InMux
    port map (
            O => \N__47336\,
            I => \N__47250\
        );

    \I__11172\ : InMux
    port map (
            O => \N__47335\,
            I => \N__47241\
        );

    \I__11171\ : InMux
    port map (
            O => \N__47334\,
            I => \N__47241\
        );

    \I__11170\ : InMux
    port map (
            O => \N__47333\,
            I => \N__47241\
        );

    \I__11169\ : InMux
    port map (
            O => \N__47332\,
            I => \N__47241\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__47329\,
            I => \N__47238\
        );

    \I__11167\ : InMux
    port map (
            O => \N__47328\,
            I => \N__47229\
        );

    \I__11166\ : InMux
    port map (
            O => \N__47327\,
            I => \N__47229\
        );

    \I__11165\ : InMux
    port map (
            O => \N__47326\,
            I => \N__47229\
        );

    \I__11164\ : InMux
    port map (
            O => \N__47325\,
            I => \N__47229\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__47322\,
            I => \N__47218\
        );

    \I__11162\ : LocalMux
    port map (
            O => \N__47311\,
            I => \N__47215\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__47308\,
            I => \N__47206\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__47299\,
            I => \N__47206\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__47292\,
            I => \N__47206\
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__47289\,
            I => \N__47206\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__47286\,
            I => \N__47188\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__47281\,
            I => \N__47188\
        );

    \I__11155\ : Span4Mux_v
    port map (
            O => \N__47278\,
            I => \N__47181\
        );

    \I__11154\ : LocalMux
    port map (
            O => \N__47265\,
            I => \N__47181\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__47258\,
            I => \N__47181\
        );

    \I__11152\ : InMux
    port map (
            O => \N__47257\,
            I => \N__47172\
        );

    \I__11151\ : InMux
    port map (
            O => \N__47256\,
            I => \N__47172\
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__47253\,
            I => \N__47169\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__47250\,
            I => \N__47160\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__47241\,
            I => \N__47160\
        );

    \I__11147\ : Span4Mux_h
    port map (
            O => \N__47238\,
            I => \N__47160\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__47229\,
            I => \N__47160\
        );

    \I__11145\ : InMux
    port map (
            O => \N__47228\,
            I => \N__47143\
        );

    \I__11144\ : InMux
    port map (
            O => \N__47227\,
            I => \N__47143\
        );

    \I__11143\ : InMux
    port map (
            O => \N__47226\,
            I => \N__47143\
        );

    \I__11142\ : InMux
    port map (
            O => \N__47225\,
            I => \N__47143\
        );

    \I__11141\ : InMux
    port map (
            O => \N__47224\,
            I => \N__47143\
        );

    \I__11140\ : InMux
    port map (
            O => \N__47223\,
            I => \N__47143\
        );

    \I__11139\ : InMux
    port map (
            O => \N__47222\,
            I => \N__47143\
        );

    \I__11138\ : InMux
    port map (
            O => \N__47221\,
            I => \N__47143\
        );

    \I__11137\ : Span4Mux_h
    port map (
            O => \N__47218\,
            I => \N__47136\
        );

    \I__11136\ : Span4Mux_v
    port map (
            O => \N__47215\,
            I => \N__47136\
        );

    \I__11135\ : Span4Mux_v
    port map (
            O => \N__47206\,
            I => \N__47136\
        );

    \I__11134\ : InMux
    port map (
            O => \N__47205\,
            I => \N__47119\
        );

    \I__11133\ : InMux
    port map (
            O => \N__47204\,
            I => \N__47119\
        );

    \I__11132\ : InMux
    port map (
            O => \N__47203\,
            I => \N__47119\
        );

    \I__11131\ : InMux
    port map (
            O => \N__47202\,
            I => \N__47119\
        );

    \I__11130\ : InMux
    port map (
            O => \N__47201\,
            I => \N__47119\
        );

    \I__11129\ : InMux
    port map (
            O => \N__47200\,
            I => \N__47119\
        );

    \I__11128\ : InMux
    port map (
            O => \N__47199\,
            I => \N__47119\
        );

    \I__11127\ : InMux
    port map (
            O => \N__47198\,
            I => \N__47119\
        );

    \I__11126\ : InMux
    port map (
            O => \N__47197\,
            I => \N__47110\
        );

    \I__11125\ : InMux
    port map (
            O => \N__47196\,
            I => \N__47110\
        );

    \I__11124\ : InMux
    port map (
            O => \N__47195\,
            I => \N__47110\
        );

    \I__11123\ : InMux
    port map (
            O => \N__47194\,
            I => \N__47110\
        );

    \I__11122\ : CascadeMux
    port map (
            O => \N__47193\,
            I => \N__47106\
        );

    \I__11121\ : Span4Mux_v
    port map (
            O => \N__47188\,
            I => \N__47100\
        );

    \I__11120\ : Span4Mux_v
    port map (
            O => \N__47181\,
            I => \N__47097\
        );

    \I__11119\ : InMux
    port map (
            O => \N__47180\,
            I => \N__47088\
        );

    \I__11118\ : InMux
    port map (
            O => \N__47179\,
            I => \N__47088\
        );

    \I__11117\ : InMux
    port map (
            O => \N__47178\,
            I => \N__47088\
        );

    \I__11116\ : InMux
    port map (
            O => \N__47177\,
            I => \N__47088\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__47172\,
            I => \N__47085\
        );

    \I__11114\ : Span4Mux_h
    port map (
            O => \N__47169\,
            I => \N__47072\
        );

    \I__11113\ : Span4Mux_v
    port map (
            O => \N__47160\,
            I => \N__47072\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__47143\,
            I => \N__47072\
        );

    \I__11111\ : Span4Mux_h
    port map (
            O => \N__47136\,
            I => \N__47072\
        );

    \I__11110\ : LocalMux
    port map (
            O => \N__47119\,
            I => \N__47072\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__47110\,
            I => \N__47072\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47109\,
            I => \N__47061\
        );

    \I__11107\ : InMux
    port map (
            O => \N__47106\,
            I => \N__47061\
        );

    \I__11106\ : InMux
    port map (
            O => \N__47105\,
            I => \N__47061\
        );

    \I__11105\ : InMux
    port map (
            O => \N__47104\,
            I => \N__47061\
        );

    \I__11104\ : InMux
    port map (
            O => \N__47103\,
            I => \N__47061\
        );

    \I__11103\ : Odrv4
    port map (
            O => \N__47100\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11102\ : Odrv4
    port map (
            O => \N__47097\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__47088\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11100\ : Odrv12
    port map (
            O => \N__47085\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11099\ : Odrv4
    port map (
            O => \N__47072\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11098\ : LocalMux
    port map (
            O => \N__47061\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11097\ : InMux
    port map (
            O => \N__47048\,
            I => \N__47043\
        );

    \I__11096\ : InMux
    port map (
            O => \N__47047\,
            I => \N__47040\
        );

    \I__11095\ : InMux
    port map (
            O => \N__47046\,
            I => \N__47037\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__47043\,
            I => \N__47034\
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__47040\,
            I => \N__47031\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__47037\,
            I => \N__47028\
        );

    \I__11091\ : Span12Mux_v
    port map (
            O => \N__47034\,
            I => \N__47024\
        );

    \I__11090\ : Span4Mux_h
    port map (
            O => \N__47031\,
            I => \N__47021\
        );

    \I__11089\ : Sp12to4
    port map (
            O => \N__47028\,
            I => \N__47018\
        );

    \I__11088\ : InMux
    port map (
            O => \N__47027\,
            I => \N__47015\
        );

    \I__11087\ : Odrv12
    port map (
            O => \N__47024\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11086\ : Odrv4
    port map (
            O => \N__47021\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11085\ : Odrv12
    port map (
            O => \N__47018\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__47015\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11083\ : CascadeMux
    port map (
            O => \N__47006\,
            I => \N__46999\
        );

    \I__11082\ : CascadeMux
    port map (
            O => \N__47005\,
            I => \N__46996\
        );

    \I__11081\ : CascadeMux
    port map (
            O => \N__47004\,
            I => \N__46993\
        );

    \I__11080\ : CascadeMux
    port map (
            O => \N__47003\,
            I => \N__46989\
        );

    \I__11079\ : InMux
    port map (
            O => \N__47002\,
            I => \N__46977\
        );

    \I__11078\ : InMux
    port map (
            O => \N__46999\,
            I => \N__46954\
        );

    \I__11077\ : InMux
    port map (
            O => \N__46996\,
            I => \N__46951\
        );

    \I__11076\ : InMux
    port map (
            O => \N__46993\,
            I => \N__46948\
        );

    \I__11075\ : InMux
    port map (
            O => \N__46992\,
            I => \N__46943\
        );

    \I__11074\ : InMux
    port map (
            O => \N__46989\,
            I => \N__46943\
        );

    \I__11073\ : InMux
    port map (
            O => \N__46988\,
            I => \N__46934\
        );

    \I__11072\ : InMux
    port map (
            O => \N__46987\,
            I => \N__46934\
        );

    \I__11071\ : InMux
    port map (
            O => \N__46986\,
            I => \N__46934\
        );

    \I__11070\ : InMux
    port map (
            O => \N__46985\,
            I => \N__46934\
        );

    \I__11069\ : InMux
    port map (
            O => \N__46984\,
            I => \N__46927\
        );

    \I__11068\ : InMux
    port map (
            O => \N__46983\,
            I => \N__46927\
        );

    \I__11067\ : InMux
    port map (
            O => \N__46982\,
            I => \N__46927\
        );

    \I__11066\ : CascadeMux
    port map (
            O => \N__46981\,
            I => \N__46923\
        );

    \I__11065\ : CascadeMux
    port map (
            O => \N__46980\,
            I => \N__46919\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__46977\,
            I => \N__46908\
        );

    \I__11063\ : InMux
    port map (
            O => \N__46976\,
            I => \N__46899\
        );

    \I__11062\ : InMux
    port map (
            O => \N__46975\,
            I => \N__46899\
        );

    \I__11061\ : InMux
    port map (
            O => \N__46974\,
            I => \N__46899\
        );

    \I__11060\ : InMux
    port map (
            O => \N__46973\,
            I => \N__46899\
        );

    \I__11059\ : InMux
    port map (
            O => \N__46972\,
            I => \N__46892\
        );

    \I__11058\ : InMux
    port map (
            O => \N__46971\,
            I => \N__46892\
        );

    \I__11057\ : InMux
    port map (
            O => \N__46970\,
            I => \N__46892\
        );

    \I__11056\ : InMux
    port map (
            O => \N__46969\,
            I => \N__46887\
        );

    \I__11055\ : InMux
    port map (
            O => \N__46968\,
            I => \N__46887\
        );

    \I__11054\ : CascadeMux
    port map (
            O => \N__46967\,
            I => \N__46868\
        );

    \I__11053\ : CascadeMux
    port map (
            O => \N__46966\,
            I => \N__46864\
        );

    \I__11052\ : CascadeMux
    port map (
            O => \N__46965\,
            I => \N__46860\
        );

    \I__11051\ : CascadeMux
    port map (
            O => \N__46964\,
            I => \N__46856\
        );

    \I__11050\ : CascadeMux
    port map (
            O => \N__46963\,
            I => \N__46852\
        );

    \I__11049\ : CascadeMux
    port map (
            O => \N__46962\,
            I => \N__46848\
        );

    \I__11048\ : CascadeMux
    port map (
            O => \N__46961\,
            I => \N__46844\
        );

    \I__11047\ : CascadeMux
    port map (
            O => \N__46960\,
            I => \N__46840\
        );

    \I__11046\ : CascadeMux
    port map (
            O => \N__46959\,
            I => \N__46836\
        );

    \I__11045\ : CascadeMux
    port map (
            O => \N__46958\,
            I => \N__46832\
        );

    \I__11044\ : CascadeMux
    port map (
            O => \N__46957\,
            I => \N__46828\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__46954\,
            I => \N__46819\
        );

    \I__11042\ : LocalMux
    port map (
            O => \N__46951\,
            I => \N__46819\
        );

    \I__11041\ : LocalMux
    port map (
            O => \N__46948\,
            I => \N__46816\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__46943\,
            I => \N__46813\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__46934\,
            I => \N__46808\
        );

    \I__11038\ : LocalMux
    port map (
            O => \N__46927\,
            I => \N__46808\
        );

    \I__11037\ : InMux
    port map (
            O => \N__46926\,
            I => \N__46789\
        );

    \I__11036\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46789\
        );

    \I__11035\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46789\
        );

    \I__11034\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46789\
        );

    \I__11033\ : InMux
    port map (
            O => \N__46918\,
            I => \N__46789\
        );

    \I__11032\ : CascadeMux
    port map (
            O => \N__46917\,
            I => \N__46785\
        );

    \I__11031\ : CascadeMux
    port map (
            O => \N__46916\,
            I => \N__46781\
        );

    \I__11030\ : CascadeMux
    port map (
            O => \N__46915\,
            I => \N__46777\
        );

    \I__11029\ : CascadeMux
    port map (
            O => \N__46914\,
            I => \N__46773\
        );

    \I__11028\ : CascadeMux
    port map (
            O => \N__46913\,
            I => \N__46769\
        );

    \I__11027\ : CascadeMux
    port map (
            O => \N__46912\,
            I => \N__46765\
        );

    \I__11026\ : CascadeMux
    port map (
            O => \N__46911\,
            I => \N__46761\
        );

    \I__11025\ : Span4Mux_v
    port map (
            O => \N__46908\,
            I => \N__46751\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__46899\,
            I => \N__46751\
        );

    \I__11023\ : LocalMux
    port map (
            O => \N__46892\,
            I => \N__46748\
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__46887\,
            I => \N__46745\
        );

    \I__11021\ : InMux
    port map (
            O => \N__46886\,
            I => \N__46742\
        );

    \I__11020\ : InMux
    port map (
            O => \N__46885\,
            I => \N__46725\
        );

    \I__11019\ : InMux
    port map (
            O => \N__46884\,
            I => \N__46725\
        );

    \I__11018\ : InMux
    port map (
            O => \N__46883\,
            I => \N__46725\
        );

    \I__11017\ : InMux
    port map (
            O => \N__46882\,
            I => \N__46725\
        );

    \I__11016\ : InMux
    port map (
            O => \N__46881\,
            I => \N__46725\
        );

    \I__11015\ : InMux
    port map (
            O => \N__46880\,
            I => \N__46725\
        );

    \I__11014\ : InMux
    port map (
            O => \N__46879\,
            I => \N__46725\
        );

    \I__11013\ : InMux
    port map (
            O => \N__46878\,
            I => \N__46725\
        );

    \I__11012\ : InMux
    port map (
            O => \N__46877\,
            I => \N__46714\
        );

    \I__11011\ : InMux
    port map (
            O => \N__46876\,
            I => \N__46714\
        );

    \I__11010\ : InMux
    port map (
            O => \N__46875\,
            I => \N__46714\
        );

    \I__11009\ : InMux
    port map (
            O => \N__46874\,
            I => \N__46714\
        );

    \I__11008\ : InMux
    port map (
            O => \N__46873\,
            I => \N__46714\
        );

    \I__11007\ : InMux
    port map (
            O => \N__46872\,
            I => \N__46697\
        );

    \I__11006\ : InMux
    port map (
            O => \N__46871\,
            I => \N__46697\
        );

    \I__11005\ : InMux
    port map (
            O => \N__46868\,
            I => \N__46697\
        );

    \I__11004\ : InMux
    port map (
            O => \N__46867\,
            I => \N__46697\
        );

    \I__11003\ : InMux
    port map (
            O => \N__46864\,
            I => \N__46697\
        );

    \I__11002\ : InMux
    port map (
            O => \N__46863\,
            I => \N__46697\
        );

    \I__11001\ : InMux
    port map (
            O => \N__46860\,
            I => \N__46697\
        );

    \I__11000\ : InMux
    port map (
            O => \N__46859\,
            I => \N__46697\
        );

    \I__10999\ : InMux
    port map (
            O => \N__46856\,
            I => \N__46680\
        );

    \I__10998\ : InMux
    port map (
            O => \N__46855\,
            I => \N__46680\
        );

    \I__10997\ : InMux
    port map (
            O => \N__46852\,
            I => \N__46680\
        );

    \I__10996\ : InMux
    port map (
            O => \N__46851\,
            I => \N__46680\
        );

    \I__10995\ : InMux
    port map (
            O => \N__46848\,
            I => \N__46680\
        );

    \I__10994\ : InMux
    port map (
            O => \N__46847\,
            I => \N__46680\
        );

    \I__10993\ : InMux
    port map (
            O => \N__46844\,
            I => \N__46680\
        );

    \I__10992\ : InMux
    port map (
            O => \N__46843\,
            I => \N__46680\
        );

    \I__10991\ : InMux
    port map (
            O => \N__46840\,
            I => \N__46663\
        );

    \I__10990\ : InMux
    port map (
            O => \N__46839\,
            I => \N__46663\
        );

    \I__10989\ : InMux
    port map (
            O => \N__46836\,
            I => \N__46663\
        );

    \I__10988\ : InMux
    port map (
            O => \N__46835\,
            I => \N__46663\
        );

    \I__10987\ : InMux
    port map (
            O => \N__46832\,
            I => \N__46663\
        );

    \I__10986\ : InMux
    port map (
            O => \N__46831\,
            I => \N__46663\
        );

    \I__10985\ : InMux
    port map (
            O => \N__46828\,
            I => \N__46663\
        );

    \I__10984\ : InMux
    port map (
            O => \N__46827\,
            I => \N__46663\
        );

    \I__10983\ : CascadeMux
    port map (
            O => \N__46826\,
            I => \N__46660\
        );

    \I__10982\ : CascadeMux
    port map (
            O => \N__46825\,
            I => \N__46656\
        );

    \I__10981\ : CascadeMux
    port map (
            O => \N__46824\,
            I => \N__46652\
        );

    \I__10980\ : Span4Mux_v
    port map (
            O => \N__46819\,
            I => \N__46645\
        );

    \I__10979\ : Span4Mux_v
    port map (
            O => \N__46816\,
            I => \N__46642\
        );

    \I__10978\ : Span4Mux_h
    port map (
            O => \N__46813\,
            I => \N__46637\
        );

    \I__10977\ : Span4Mux_h
    port map (
            O => \N__46808\,
            I => \N__46637\
        );

    \I__10976\ : CascadeMux
    port map (
            O => \N__46807\,
            I => \N__46634\
        );

    \I__10975\ : CascadeMux
    port map (
            O => \N__46806\,
            I => \N__46629\
        );

    \I__10974\ : CascadeMux
    port map (
            O => \N__46805\,
            I => \N__46625\
        );

    \I__10973\ : CascadeMux
    port map (
            O => \N__46804\,
            I => \N__46622\
        );

    \I__10972\ : CascadeMux
    port map (
            O => \N__46803\,
            I => \N__46619\
        );

    \I__10971\ : CascadeMux
    port map (
            O => \N__46802\,
            I => \N__46614\
        );

    \I__10970\ : CascadeMux
    port map (
            O => \N__46801\,
            I => \N__46610\
        );

    \I__10969\ : CascadeMux
    port map (
            O => \N__46800\,
            I => \N__46607\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__46789\,
            I => \N__46602\
        );

    \I__10967\ : InMux
    port map (
            O => \N__46788\,
            I => \N__46587\
        );

    \I__10966\ : InMux
    port map (
            O => \N__46785\,
            I => \N__46587\
        );

    \I__10965\ : InMux
    port map (
            O => \N__46784\,
            I => \N__46587\
        );

    \I__10964\ : InMux
    port map (
            O => \N__46781\,
            I => \N__46587\
        );

    \I__10963\ : InMux
    port map (
            O => \N__46780\,
            I => \N__46587\
        );

    \I__10962\ : InMux
    port map (
            O => \N__46777\,
            I => \N__46587\
        );

    \I__10961\ : InMux
    port map (
            O => \N__46776\,
            I => \N__46587\
        );

    \I__10960\ : InMux
    port map (
            O => \N__46773\,
            I => \N__46570\
        );

    \I__10959\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46570\
        );

    \I__10958\ : InMux
    port map (
            O => \N__46769\,
            I => \N__46570\
        );

    \I__10957\ : InMux
    port map (
            O => \N__46768\,
            I => \N__46570\
        );

    \I__10956\ : InMux
    port map (
            O => \N__46765\,
            I => \N__46570\
        );

    \I__10955\ : InMux
    port map (
            O => \N__46764\,
            I => \N__46570\
        );

    \I__10954\ : InMux
    port map (
            O => \N__46761\,
            I => \N__46570\
        );

    \I__10953\ : InMux
    port map (
            O => \N__46760\,
            I => \N__46570\
        );

    \I__10952\ : CascadeMux
    port map (
            O => \N__46759\,
            I => \N__46567\
        );

    \I__10951\ : CascadeMux
    port map (
            O => \N__46758\,
            I => \N__46563\
        );

    \I__10950\ : CascadeMux
    port map (
            O => \N__46757\,
            I => \N__46559\
        );

    \I__10949\ : CascadeMux
    port map (
            O => \N__46756\,
            I => \N__46555\
        );

    \I__10948\ : Span4Mux_h
    port map (
            O => \N__46751\,
            I => \N__46543\
        );

    \I__10947\ : Span4Mux_h
    port map (
            O => \N__46748\,
            I => \N__46543\
        );

    \I__10946\ : Span4Mux_v
    port map (
            O => \N__46745\,
            I => \N__46543\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__46742\,
            I => \N__46543\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__46725\,
            I => \N__46543\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__46714\,
            I => \N__46534\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__46697\,
            I => \N__46534\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__46680\,
            I => \N__46534\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__46663\,
            I => \N__46534\
        );

    \I__10939\ : InMux
    port map (
            O => \N__46660\,
            I => \N__46521\
        );

    \I__10938\ : InMux
    port map (
            O => \N__46659\,
            I => \N__46521\
        );

    \I__10937\ : InMux
    port map (
            O => \N__46656\,
            I => \N__46521\
        );

    \I__10936\ : InMux
    port map (
            O => \N__46655\,
            I => \N__46521\
        );

    \I__10935\ : InMux
    port map (
            O => \N__46652\,
            I => \N__46521\
        );

    \I__10934\ : InMux
    port map (
            O => \N__46651\,
            I => \N__46521\
        );

    \I__10933\ : CascadeMux
    port map (
            O => \N__46650\,
            I => \N__46518\
        );

    \I__10932\ : CascadeMux
    port map (
            O => \N__46649\,
            I => \N__46514\
        );

    \I__10931\ : CascadeMux
    port map (
            O => \N__46648\,
            I => \N__46510\
        );

    \I__10930\ : Span4Mux_v
    port map (
            O => \N__46645\,
            I => \N__46504\
        );

    \I__10929\ : Span4Mux_v
    port map (
            O => \N__46642\,
            I => \N__46504\
        );

    \I__10928\ : Span4Mux_v
    port map (
            O => \N__46637\,
            I => \N__46501\
        );

    \I__10927\ : InMux
    port map (
            O => \N__46634\,
            I => \N__46490\
        );

    \I__10926\ : InMux
    port map (
            O => \N__46633\,
            I => \N__46490\
        );

    \I__10925\ : InMux
    port map (
            O => \N__46632\,
            I => \N__46490\
        );

    \I__10924\ : InMux
    port map (
            O => \N__46629\,
            I => \N__46490\
        );

    \I__10923\ : InMux
    port map (
            O => \N__46628\,
            I => \N__46490\
        );

    \I__10922\ : InMux
    port map (
            O => \N__46625\,
            I => \N__46483\
        );

    \I__10921\ : InMux
    port map (
            O => \N__46622\,
            I => \N__46483\
        );

    \I__10920\ : InMux
    port map (
            O => \N__46619\,
            I => \N__46483\
        );

    \I__10919\ : InMux
    port map (
            O => \N__46618\,
            I => \N__46474\
        );

    \I__10918\ : InMux
    port map (
            O => \N__46617\,
            I => \N__46474\
        );

    \I__10917\ : InMux
    port map (
            O => \N__46614\,
            I => \N__46474\
        );

    \I__10916\ : InMux
    port map (
            O => \N__46613\,
            I => \N__46474\
        );

    \I__10915\ : InMux
    port map (
            O => \N__46610\,
            I => \N__46469\
        );

    \I__10914\ : InMux
    port map (
            O => \N__46607\,
            I => \N__46469\
        );

    \I__10913\ : InMux
    port map (
            O => \N__46606\,
            I => \N__46464\
        );

    \I__10912\ : InMux
    port map (
            O => \N__46605\,
            I => \N__46464\
        );

    \I__10911\ : Span4Mux_h
    port map (
            O => \N__46602\,
            I => \N__46457\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__46587\,
            I => \N__46457\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__46570\,
            I => \N__46457\
        );

    \I__10908\ : InMux
    port map (
            O => \N__46567\,
            I => \N__46440\
        );

    \I__10907\ : InMux
    port map (
            O => \N__46566\,
            I => \N__46440\
        );

    \I__10906\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46440\
        );

    \I__10905\ : InMux
    port map (
            O => \N__46562\,
            I => \N__46440\
        );

    \I__10904\ : InMux
    port map (
            O => \N__46559\,
            I => \N__46440\
        );

    \I__10903\ : InMux
    port map (
            O => \N__46558\,
            I => \N__46440\
        );

    \I__10902\ : InMux
    port map (
            O => \N__46555\,
            I => \N__46440\
        );

    \I__10901\ : InMux
    port map (
            O => \N__46554\,
            I => \N__46440\
        );

    \I__10900\ : Span4Mux_v
    port map (
            O => \N__46543\,
            I => \N__46433\
        );

    \I__10899\ : Span4Mux_v
    port map (
            O => \N__46534\,
            I => \N__46433\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__46521\,
            I => \N__46433\
        );

    \I__10897\ : InMux
    port map (
            O => \N__46518\,
            I => \N__46420\
        );

    \I__10896\ : InMux
    port map (
            O => \N__46517\,
            I => \N__46420\
        );

    \I__10895\ : InMux
    port map (
            O => \N__46514\,
            I => \N__46420\
        );

    \I__10894\ : InMux
    port map (
            O => \N__46513\,
            I => \N__46420\
        );

    \I__10893\ : InMux
    port map (
            O => \N__46510\,
            I => \N__46420\
        );

    \I__10892\ : InMux
    port map (
            O => \N__46509\,
            I => \N__46420\
        );

    \I__10891\ : Odrv4
    port map (
            O => \N__46504\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10890\ : Odrv4
    port map (
            O => \N__46501\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__46490\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__46483\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__46474\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__46469\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__46464\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10884\ : Odrv4
    port map (
            O => \N__46457\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__46440\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10882\ : Odrv4
    port map (
            O => \N__46433\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__46420\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10880\ : CascadeMux
    port map (
            O => \N__46397\,
            I => \N__46394\
        );

    \I__10879\ : InMux
    port map (
            O => \N__46394\,
            I => \N__46390\
        );

    \I__10878\ : InMux
    port map (
            O => \N__46393\,
            I => \N__46386\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__46390\,
            I => \N__46383\
        );

    \I__10876\ : InMux
    port map (
            O => \N__46389\,
            I => \N__46380\
        );

    \I__10875\ : LocalMux
    port map (
            O => \N__46386\,
            I => \N__46377\
        );

    \I__10874\ : Span4Mux_h
    port map (
            O => \N__46383\,
            I => \N__46374\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__46380\,
            I => \N__46371\
        );

    \I__10872\ : Odrv12
    port map (
            O => \N__46377\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__10871\ : Odrv4
    port map (
            O => \N__46374\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__10870\ : Odrv12
    port map (
            O => \N__46371\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__10869\ : InMux
    port map (
            O => \N__46364\,
            I => \N__46361\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__46361\,
            I => \N__46358\
        );

    \I__10867\ : Odrv4
    port map (
            O => \N__46358\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__10866\ : InMux
    port map (
            O => \N__46355\,
            I => \N__46352\
        );

    \I__10865\ : LocalMux
    port map (
            O => \N__46352\,
            I => \N__46347\
        );

    \I__10864\ : InMux
    port map (
            O => \N__46351\,
            I => \N__46344\
        );

    \I__10863\ : InMux
    port map (
            O => \N__46350\,
            I => \N__46341\
        );

    \I__10862\ : Span4Mux_h
    port map (
            O => \N__46347\,
            I => \N__46338\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__46344\,
            I => \N__46335\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__46341\,
            I => \N__46332\
        );

    \I__10859\ : Span4Mux_v
    port map (
            O => \N__46338\,
            I => \N__46329\
        );

    \I__10858\ : Span4Mux_h
    port map (
            O => \N__46335\,
            I => \N__46326\
        );

    \I__10857\ : Span4Mux_h
    port map (
            O => \N__46332\,
            I => \N__46323\
        );

    \I__10856\ : Span4Mux_v
    port map (
            O => \N__46329\,
            I => \N__46320\
        );

    \I__10855\ : Sp12to4
    port map (
            O => \N__46326\,
            I => \N__46317\
        );

    \I__10854\ : Span4Mux_v
    port map (
            O => \N__46323\,
            I => \N__46314\
        );

    \I__10853\ : Span4Mux_v
    port map (
            O => \N__46320\,
            I => \N__46311\
        );

    \I__10852\ : Span12Mux_v
    port map (
            O => \N__46317\,
            I => \N__46308\
        );

    \I__10851\ : Sp12to4
    port map (
            O => \N__46314\,
            I => \N__46305\
        );

    \I__10850\ : Span4Mux_v
    port map (
            O => \N__46311\,
            I => \N__46302\
        );

    \I__10849\ : Span12Mux_v
    port map (
            O => \N__46308\,
            I => \N__46299\
        );

    \I__10848\ : Span12Mux_v
    port map (
            O => \N__46305\,
            I => \N__46296\
        );

    \I__10847\ : Span4Mux_v
    port map (
            O => \N__46302\,
            I => \N__46293\
        );

    \I__10846\ : Odrv12
    port map (
            O => \N__46299\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__10845\ : Odrv12
    port map (
            O => \N__46296\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__10844\ : Odrv4
    port map (
            O => \N__46293\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__10843\ : InMux
    port map (
            O => \N__46286\,
            I => \N__46282\
        );

    \I__10842\ : InMux
    port map (
            O => \N__46285\,
            I => \N__46279\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__46282\,
            I => \N__46274\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__46279\,
            I => \N__46274\
        );

    \I__10839\ : Span12Mux_v
    port map (
            O => \N__46274\,
            I => \N__46269\
        );

    \I__10838\ : InMux
    port map (
            O => \N__46273\,
            I => \N__46264\
        );

    \I__10837\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46264\
        );

    \I__10836\ : Span12Mux_v
    port map (
            O => \N__46269\,
            I => \N__46261\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__46264\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__10834\ : Odrv12
    port map (
            O => \N__46261\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__10833\ : ClkMux
    port map (
            O => \N__46256\,
            I => \N__46253\
        );

    \I__10832\ : GlobalMux
    port map (
            O => \N__46253\,
            I => \N__46250\
        );

    \I__10831\ : gio2CtrlBuf
    port map (
            O => \N__46250\,
            I => delay_tr_input_c_g
        );

    \I__10830\ : CascadeMux
    port map (
            O => \N__46247\,
            I => \N__46244\
        );

    \I__10829\ : InMux
    port map (
            O => \N__46244\,
            I => \N__46240\
        );

    \I__10828\ : InMux
    port map (
            O => \N__46243\,
            I => \N__46237\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__46240\,
            I => \N__46234\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__46237\,
            I => \N__46230\
        );

    \I__10825\ : Span4Mux_v
    port map (
            O => \N__46234\,
            I => \N__46225\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46233\,
            I => \N__46222\
        );

    \I__10823\ : Span4Mux_h
    port map (
            O => \N__46230\,
            I => \N__46218\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46229\,
            I => \N__46215\
        );

    \I__10821\ : InMux
    port map (
            O => \N__46228\,
            I => \N__46212\
        );

    \I__10820\ : Span4Mux_h
    port map (
            O => \N__46225\,
            I => \N__46207\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__46222\,
            I => \N__46207\
        );

    \I__10818\ : CascadeMux
    port map (
            O => \N__46221\,
            I => \N__46204\
        );

    \I__10817\ : Span4Mux_h
    port map (
            O => \N__46218\,
            I => \N__46201\
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__46215\,
            I => \N__46196\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__46212\,
            I => \N__46196\
        );

    \I__10814\ : Span4Mux_v
    port map (
            O => \N__46207\,
            I => \N__46193\
        );

    \I__10813\ : InMux
    port map (
            O => \N__46204\,
            I => \N__46190\
        );

    \I__10812\ : Span4Mux_v
    port map (
            O => \N__46201\,
            I => \N__46187\
        );

    \I__10811\ : Span4Mux_v
    port map (
            O => \N__46196\,
            I => \N__46182\
        );

    \I__10810\ : Span4Mux_v
    port map (
            O => \N__46193\,
            I => \N__46182\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__46190\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__10808\ : Odrv4
    port map (
            O => \N__46187\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__10807\ : Odrv4
    port map (
            O => \N__46182\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__10806\ : InMux
    port map (
            O => \N__46175\,
            I => \N__46172\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46172\,
            I => \N__46169\
        );

    \I__10804\ : Span4Mux_v
    port map (
            O => \N__46169\,
            I => \N__46165\
        );

    \I__10803\ : InMux
    port map (
            O => \N__46168\,
            I => \N__46162\
        );

    \I__10802\ : Span4Mux_h
    port map (
            O => \N__46165\,
            I => \N__46159\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__46162\,
            I => \N__46156\
        );

    \I__10800\ : Span4Mux_v
    port map (
            O => \N__46159\,
            I => \N__46153\
        );

    \I__10799\ : Span4Mux_h
    port map (
            O => \N__46156\,
            I => \N__46148\
        );

    \I__10798\ : Span4Mux_v
    port map (
            O => \N__46153\,
            I => \N__46145\
        );

    \I__10797\ : InMux
    port map (
            O => \N__46152\,
            I => \N__46140\
        );

    \I__10796\ : InMux
    port map (
            O => \N__46151\,
            I => \N__46140\
        );

    \I__10795\ : Odrv4
    port map (
            O => \N__46148\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__10794\ : Odrv4
    port map (
            O => \N__46145\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__46140\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__10792\ : IoInMux
    port map (
            O => \N__46133\,
            I => \N__46130\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__46130\,
            I => \N__46126\
        );

    \I__10790\ : InMux
    port map (
            O => \N__46129\,
            I => \N__46123\
        );

    \I__10789\ : Odrv12
    port map (
            O => \N__46126\,
            I => \T23_c\
        );

    \I__10788\ : LocalMux
    port map (
            O => \N__46123\,
            I => \T23_c\
        );

    \I__10787\ : ClkMux
    port map (
            O => \N__46118\,
            I => \N__45731\
        );

    \I__10786\ : ClkMux
    port map (
            O => \N__46117\,
            I => \N__45731\
        );

    \I__10785\ : ClkMux
    port map (
            O => \N__46116\,
            I => \N__45731\
        );

    \I__10784\ : ClkMux
    port map (
            O => \N__46115\,
            I => \N__45731\
        );

    \I__10783\ : ClkMux
    port map (
            O => \N__46114\,
            I => \N__45731\
        );

    \I__10782\ : ClkMux
    port map (
            O => \N__46113\,
            I => \N__45731\
        );

    \I__10781\ : ClkMux
    port map (
            O => \N__46112\,
            I => \N__45731\
        );

    \I__10780\ : ClkMux
    port map (
            O => \N__46111\,
            I => \N__45731\
        );

    \I__10779\ : ClkMux
    port map (
            O => \N__46110\,
            I => \N__45731\
        );

    \I__10778\ : ClkMux
    port map (
            O => \N__46109\,
            I => \N__45731\
        );

    \I__10777\ : ClkMux
    port map (
            O => \N__46108\,
            I => \N__45731\
        );

    \I__10776\ : ClkMux
    port map (
            O => \N__46107\,
            I => \N__45731\
        );

    \I__10775\ : ClkMux
    port map (
            O => \N__46106\,
            I => \N__45731\
        );

    \I__10774\ : ClkMux
    port map (
            O => \N__46105\,
            I => \N__45731\
        );

    \I__10773\ : ClkMux
    port map (
            O => \N__46104\,
            I => \N__45731\
        );

    \I__10772\ : ClkMux
    port map (
            O => \N__46103\,
            I => \N__45731\
        );

    \I__10771\ : ClkMux
    port map (
            O => \N__46102\,
            I => \N__45731\
        );

    \I__10770\ : ClkMux
    port map (
            O => \N__46101\,
            I => \N__45731\
        );

    \I__10769\ : ClkMux
    port map (
            O => \N__46100\,
            I => \N__45731\
        );

    \I__10768\ : ClkMux
    port map (
            O => \N__46099\,
            I => \N__45731\
        );

    \I__10767\ : ClkMux
    port map (
            O => \N__46098\,
            I => \N__45731\
        );

    \I__10766\ : ClkMux
    port map (
            O => \N__46097\,
            I => \N__45731\
        );

    \I__10765\ : ClkMux
    port map (
            O => \N__46096\,
            I => \N__45731\
        );

    \I__10764\ : ClkMux
    port map (
            O => \N__46095\,
            I => \N__45731\
        );

    \I__10763\ : ClkMux
    port map (
            O => \N__46094\,
            I => \N__45731\
        );

    \I__10762\ : ClkMux
    port map (
            O => \N__46093\,
            I => \N__45731\
        );

    \I__10761\ : ClkMux
    port map (
            O => \N__46092\,
            I => \N__45731\
        );

    \I__10760\ : ClkMux
    port map (
            O => \N__46091\,
            I => \N__45731\
        );

    \I__10759\ : ClkMux
    port map (
            O => \N__46090\,
            I => \N__45731\
        );

    \I__10758\ : ClkMux
    port map (
            O => \N__46089\,
            I => \N__45731\
        );

    \I__10757\ : ClkMux
    port map (
            O => \N__46088\,
            I => \N__45731\
        );

    \I__10756\ : ClkMux
    port map (
            O => \N__46087\,
            I => \N__45731\
        );

    \I__10755\ : ClkMux
    port map (
            O => \N__46086\,
            I => \N__45731\
        );

    \I__10754\ : ClkMux
    port map (
            O => \N__46085\,
            I => \N__45731\
        );

    \I__10753\ : ClkMux
    port map (
            O => \N__46084\,
            I => \N__45731\
        );

    \I__10752\ : ClkMux
    port map (
            O => \N__46083\,
            I => \N__45731\
        );

    \I__10751\ : ClkMux
    port map (
            O => \N__46082\,
            I => \N__45731\
        );

    \I__10750\ : ClkMux
    port map (
            O => \N__46081\,
            I => \N__45731\
        );

    \I__10749\ : ClkMux
    port map (
            O => \N__46080\,
            I => \N__45731\
        );

    \I__10748\ : ClkMux
    port map (
            O => \N__46079\,
            I => \N__45731\
        );

    \I__10747\ : ClkMux
    port map (
            O => \N__46078\,
            I => \N__45731\
        );

    \I__10746\ : ClkMux
    port map (
            O => \N__46077\,
            I => \N__45731\
        );

    \I__10745\ : ClkMux
    port map (
            O => \N__46076\,
            I => \N__45731\
        );

    \I__10744\ : ClkMux
    port map (
            O => \N__46075\,
            I => \N__45731\
        );

    \I__10743\ : ClkMux
    port map (
            O => \N__46074\,
            I => \N__45731\
        );

    \I__10742\ : ClkMux
    port map (
            O => \N__46073\,
            I => \N__45731\
        );

    \I__10741\ : ClkMux
    port map (
            O => \N__46072\,
            I => \N__45731\
        );

    \I__10740\ : ClkMux
    port map (
            O => \N__46071\,
            I => \N__45731\
        );

    \I__10739\ : ClkMux
    port map (
            O => \N__46070\,
            I => \N__45731\
        );

    \I__10738\ : ClkMux
    port map (
            O => \N__46069\,
            I => \N__45731\
        );

    \I__10737\ : ClkMux
    port map (
            O => \N__46068\,
            I => \N__45731\
        );

    \I__10736\ : ClkMux
    port map (
            O => \N__46067\,
            I => \N__45731\
        );

    \I__10735\ : ClkMux
    port map (
            O => \N__46066\,
            I => \N__45731\
        );

    \I__10734\ : ClkMux
    port map (
            O => \N__46065\,
            I => \N__45731\
        );

    \I__10733\ : ClkMux
    port map (
            O => \N__46064\,
            I => \N__45731\
        );

    \I__10732\ : ClkMux
    port map (
            O => \N__46063\,
            I => \N__45731\
        );

    \I__10731\ : ClkMux
    port map (
            O => \N__46062\,
            I => \N__45731\
        );

    \I__10730\ : ClkMux
    port map (
            O => \N__46061\,
            I => \N__45731\
        );

    \I__10729\ : ClkMux
    port map (
            O => \N__46060\,
            I => \N__45731\
        );

    \I__10728\ : ClkMux
    port map (
            O => \N__46059\,
            I => \N__45731\
        );

    \I__10727\ : ClkMux
    port map (
            O => \N__46058\,
            I => \N__45731\
        );

    \I__10726\ : ClkMux
    port map (
            O => \N__46057\,
            I => \N__45731\
        );

    \I__10725\ : ClkMux
    port map (
            O => \N__46056\,
            I => \N__45731\
        );

    \I__10724\ : ClkMux
    port map (
            O => \N__46055\,
            I => \N__45731\
        );

    \I__10723\ : ClkMux
    port map (
            O => \N__46054\,
            I => \N__45731\
        );

    \I__10722\ : ClkMux
    port map (
            O => \N__46053\,
            I => \N__45731\
        );

    \I__10721\ : ClkMux
    port map (
            O => \N__46052\,
            I => \N__45731\
        );

    \I__10720\ : ClkMux
    port map (
            O => \N__46051\,
            I => \N__45731\
        );

    \I__10719\ : ClkMux
    port map (
            O => \N__46050\,
            I => \N__45731\
        );

    \I__10718\ : ClkMux
    port map (
            O => \N__46049\,
            I => \N__45731\
        );

    \I__10717\ : ClkMux
    port map (
            O => \N__46048\,
            I => \N__45731\
        );

    \I__10716\ : ClkMux
    port map (
            O => \N__46047\,
            I => \N__45731\
        );

    \I__10715\ : ClkMux
    port map (
            O => \N__46046\,
            I => \N__45731\
        );

    \I__10714\ : ClkMux
    port map (
            O => \N__46045\,
            I => \N__45731\
        );

    \I__10713\ : ClkMux
    port map (
            O => \N__46044\,
            I => \N__45731\
        );

    \I__10712\ : ClkMux
    port map (
            O => \N__46043\,
            I => \N__45731\
        );

    \I__10711\ : ClkMux
    port map (
            O => \N__46042\,
            I => \N__45731\
        );

    \I__10710\ : ClkMux
    port map (
            O => \N__46041\,
            I => \N__45731\
        );

    \I__10709\ : ClkMux
    port map (
            O => \N__46040\,
            I => \N__45731\
        );

    \I__10708\ : ClkMux
    port map (
            O => \N__46039\,
            I => \N__45731\
        );

    \I__10707\ : ClkMux
    port map (
            O => \N__46038\,
            I => \N__45731\
        );

    \I__10706\ : ClkMux
    port map (
            O => \N__46037\,
            I => \N__45731\
        );

    \I__10705\ : ClkMux
    port map (
            O => \N__46036\,
            I => \N__45731\
        );

    \I__10704\ : ClkMux
    port map (
            O => \N__46035\,
            I => \N__45731\
        );

    \I__10703\ : ClkMux
    port map (
            O => \N__46034\,
            I => \N__45731\
        );

    \I__10702\ : ClkMux
    port map (
            O => \N__46033\,
            I => \N__45731\
        );

    \I__10701\ : ClkMux
    port map (
            O => \N__46032\,
            I => \N__45731\
        );

    \I__10700\ : ClkMux
    port map (
            O => \N__46031\,
            I => \N__45731\
        );

    \I__10699\ : ClkMux
    port map (
            O => \N__46030\,
            I => \N__45731\
        );

    \I__10698\ : ClkMux
    port map (
            O => \N__46029\,
            I => \N__45731\
        );

    \I__10697\ : ClkMux
    port map (
            O => \N__46028\,
            I => \N__45731\
        );

    \I__10696\ : ClkMux
    port map (
            O => \N__46027\,
            I => \N__45731\
        );

    \I__10695\ : ClkMux
    port map (
            O => \N__46026\,
            I => \N__45731\
        );

    \I__10694\ : ClkMux
    port map (
            O => \N__46025\,
            I => \N__45731\
        );

    \I__10693\ : ClkMux
    port map (
            O => \N__46024\,
            I => \N__45731\
        );

    \I__10692\ : ClkMux
    port map (
            O => \N__46023\,
            I => \N__45731\
        );

    \I__10691\ : ClkMux
    port map (
            O => \N__46022\,
            I => \N__45731\
        );

    \I__10690\ : ClkMux
    port map (
            O => \N__46021\,
            I => \N__45731\
        );

    \I__10689\ : ClkMux
    port map (
            O => \N__46020\,
            I => \N__45731\
        );

    \I__10688\ : ClkMux
    port map (
            O => \N__46019\,
            I => \N__45731\
        );

    \I__10687\ : ClkMux
    port map (
            O => \N__46018\,
            I => \N__45731\
        );

    \I__10686\ : ClkMux
    port map (
            O => \N__46017\,
            I => \N__45731\
        );

    \I__10685\ : ClkMux
    port map (
            O => \N__46016\,
            I => \N__45731\
        );

    \I__10684\ : ClkMux
    port map (
            O => \N__46015\,
            I => \N__45731\
        );

    \I__10683\ : ClkMux
    port map (
            O => \N__46014\,
            I => \N__45731\
        );

    \I__10682\ : ClkMux
    port map (
            O => \N__46013\,
            I => \N__45731\
        );

    \I__10681\ : ClkMux
    port map (
            O => \N__46012\,
            I => \N__45731\
        );

    \I__10680\ : ClkMux
    port map (
            O => \N__46011\,
            I => \N__45731\
        );

    \I__10679\ : ClkMux
    port map (
            O => \N__46010\,
            I => \N__45731\
        );

    \I__10678\ : ClkMux
    port map (
            O => \N__46009\,
            I => \N__45731\
        );

    \I__10677\ : ClkMux
    port map (
            O => \N__46008\,
            I => \N__45731\
        );

    \I__10676\ : ClkMux
    port map (
            O => \N__46007\,
            I => \N__45731\
        );

    \I__10675\ : ClkMux
    port map (
            O => \N__46006\,
            I => \N__45731\
        );

    \I__10674\ : ClkMux
    port map (
            O => \N__46005\,
            I => \N__45731\
        );

    \I__10673\ : ClkMux
    port map (
            O => \N__46004\,
            I => \N__45731\
        );

    \I__10672\ : ClkMux
    port map (
            O => \N__46003\,
            I => \N__45731\
        );

    \I__10671\ : ClkMux
    port map (
            O => \N__46002\,
            I => \N__45731\
        );

    \I__10670\ : ClkMux
    port map (
            O => \N__46001\,
            I => \N__45731\
        );

    \I__10669\ : ClkMux
    port map (
            O => \N__46000\,
            I => \N__45731\
        );

    \I__10668\ : ClkMux
    port map (
            O => \N__45999\,
            I => \N__45731\
        );

    \I__10667\ : ClkMux
    port map (
            O => \N__45998\,
            I => \N__45731\
        );

    \I__10666\ : ClkMux
    port map (
            O => \N__45997\,
            I => \N__45731\
        );

    \I__10665\ : ClkMux
    port map (
            O => \N__45996\,
            I => \N__45731\
        );

    \I__10664\ : ClkMux
    port map (
            O => \N__45995\,
            I => \N__45731\
        );

    \I__10663\ : ClkMux
    port map (
            O => \N__45994\,
            I => \N__45731\
        );

    \I__10662\ : ClkMux
    port map (
            O => \N__45993\,
            I => \N__45731\
        );

    \I__10661\ : ClkMux
    port map (
            O => \N__45992\,
            I => \N__45731\
        );

    \I__10660\ : ClkMux
    port map (
            O => \N__45991\,
            I => \N__45731\
        );

    \I__10659\ : ClkMux
    port map (
            O => \N__45990\,
            I => \N__45731\
        );

    \I__10658\ : GlobalMux
    port map (
            O => \N__45731\,
            I => clk_100mhz_0
        );

    \I__10657\ : InMux
    port map (
            O => \N__45728\,
            I => \N__45711\
        );

    \I__10656\ : InMux
    port map (
            O => \N__45727\,
            I => \N__45708\
        );

    \I__10655\ : InMux
    port map (
            O => \N__45726\,
            I => \N__45705\
        );

    \I__10654\ : InMux
    port map (
            O => \N__45725\,
            I => \N__45702\
        );

    \I__10653\ : InMux
    port map (
            O => \N__45724\,
            I => \N__45699\
        );

    \I__10652\ : InMux
    port map (
            O => \N__45723\,
            I => \N__45694\
        );

    \I__10651\ : InMux
    port map (
            O => \N__45722\,
            I => \N__45694\
        );

    \I__10650\ : InMux
    port map (
            O => \N__45721\,
            I => \N__45691\
        );

    \I__10649\ : InMux
    port map (
            O => \N__45720\,
            I => \N__45686\
        );

    \I__10648\ : InMux
    port map (
            O => \N__45719\,
            I => \N__45686\
        );

    \I__10647\ : InMux
    port map (
            O => \N__45718\,
            I => \N__45683\
        );

    \I__10646\ : InMux
    port map (
            O => \N__45717\,
            I => \N__45678\
        );

    \I__10645\ : InMux
    port map (
            O => \N__45716\,
            I => \N__45678\
        );

    \I__10644\ : InMux
    port map (
            O => \N__45715\,
            I => \N__45675\
        );

    \I__10643\ : InMux
    port map (
            O => \N__45714\,
            I => \N__45672\
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__45711\,
            I => \N__45669\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__45708\,
            I => \N__45666\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__45705\,
            I => \N__45663\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__45702\,
            I => \N__45659\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__45699\,
            I => \N__45646\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__45694\,
            I => \N__45643\
        );

    \I__10636\ : LocalMux
    port map (
            O => \N__45691\,
            I => \N__45627\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__45686\,
            I => \N__45616\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__45683\,
            I => \N__45613\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__45678\,
            I => \N__45523\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__45675\,
            I => \N__45520\
        );

    \I__10631\ : LocalMux
    port map (
            O => \N__45672\,
            I => \N__45516\
        );

    \I__10630\ : Glb2LocalMux
    port map (
            O => \N__45669\,
            I => \N__45245\
        );

    \I__10629\ : Glb2LocalMux
    port map (
            O => \N__45666\,
            I => \N__45245\
        );

    \I__10628\ : Glb2LocalMux
    port map (
            O => \N__45663\,
            I => \N__45245\
        );

    \I__10627\ : SRMux
    port map (
            O => \N__45662\,
            I => \N__45245\
        );

    \I__10626\ : Glb2LocalMux
    port map (
            O => \N__45659\,
            I => \N__45245\
        );

    \I__10625\ : SRMux
    port map (
            O => \N__45658\,
            I => \N__45245\
        );

    \I__10624\ : SRMux
    port map (
            O => \N__45657\,
            I => \N__45245\
        );

    \I__10623\ : SRMux
    port map (
            O => \N__45656\,
            I => \N__45245\
        );

    \I__10622\ : SRMux
    port map (
            O => \N__45655\,
            I => \N__45245\
        );

    \I__10621\ : SRMux
    port map (
            O => \N__45654\,
            I => \N__45245\
        );

    \I__10620\ : SRMux
    port map (
            O => \N__45653\,
            I => \N__45245\
        );

    \I__10619\ : SRMux
    port map (
            O => \N__45652\,
            I => \N__45245\
        );

    \I__10618\ : SRMux
    port map (
            O => \N__45651\,
            I => \N__45245\
        );

    \I__10617\ : SRMux
    port map (
            O => \N__45650\,
            I => \N__45245\
        );

    \I__10616\ : SRMux
    port map (
            O => \N__45649\,
            I => \N__45245\
        );

    \I__10615\ : Glb2LocalMux
    port map (
            O => \N__45646\,
            I => \N__45245\
        );

    \I__10614\ : Glb2LocalMux
    port map (
            O => \N__45643\,
            I => \N__45245\
        );

    \I__10613\ : SRMux
    port map (
            O => \N__45642\,
            I => \N__45245\
        );

    \I__10612\ : SRMux
    port map (
            O => \N__45641\,
            I => \N__45245\
        );

    \I__10611\ : SRMux
    port map (
            O => \N__45640\,
            I => \N__45245\
        );

    \I__10610\ : SRMux
    port map (
            O => \N__45639\,
            I => \N__45245\
        );

    \I__10609\ : SRMux
    port map (
            O => \N__45638\,
            I => \N__45245\
        );

    \I__10608\ : SRMux
    port map (
            O => \N__45637\,
            I => \N__45245\
        );

    \I__10607\ : SRMux
    port map (
            O => \N__45636\,
            I => \N__45245\
        );

    \I__10606\ : SRMux
    port map (
            O => \N__45635\,
            I => \N__45245\
        );

    \I__10605\ : SRMux
    port map (
            O => \N__45634\,
            I => \N__45245\
        );

    \I__10604\ : SRMux
    port map (
            O => \N__45633\,
            I => \N__45245\
        );

    \I__10603\ : SRMux
    port map (
            O => \N__45632\,
            I => \N__45245\
        );

    \I__10602\ : SRMux
    port map (
            O => \N__45631\,
            I => \N__45245\
        );

    \I__10601\ : SRMux
    port map (
            O => \N__45630\,
            I => \N__45245\
        );

    \I__10600\ : Glb2LocalMux
    port map (
            O => \N__45627\,
            I => \N__45245\
        );

    \I__10599\ : SRMux
    port map (
            O => \N__45626\,
            I => \N__45245\
        );

    \I__10598\ : SRMux
    port map (
            O => \N__45625\,
            I => \N__45245\
        );

    \I__10597\ : SRMux
    port map (
            O => \N__45624\,
            I => \N__45245\
        );

    \I__10596\ : SRMux
    port map (
            O => \N__45623\,
            I => \N__45245\
        );

    \I__10595\ : SRMux
    port map (
            O => \N__45622\,
            I => \N__45245\
        );

    \I__10594\ : SRMux
    port map (
            O => \N__45621\,
            I => \N__45245\
        );

    \I__10593\ : SRMux
    port map (
            O => \N__45620\,
            I => \N__45245\
        );

    \I__10592\ : SRMux
    port map (
            O => \N__45619\,
            I => \N__45245\
        );

    \I__10591\ : Glb2LocalMux
    port map (
            O => \N__45616\,
            I => \N__45245\
        );

    \I__10590\ : Glb2LocalMux
    port map (
            O => \N__45613\,
            I => \N__45245\
        );

    \I__10589\ : SRMux
    port map (
            O => \N__45612\,
            I => \N__45245\
        );

    \I__10588\ : SRMux
    port map (
            O => \N__45611\,
            I => \N__45245\
        );

    \I__10587\ : SRMux
    port map (
            O => \N__45610\,
            I => \N__45245\
        );

    \I__10586\ : SRMux
    port map (
            O => \N__45609\,
            I => \N__45245\
        );

    \I__10585\ : SRMux
    port map (
            O => \N__45608\,
            I => \N__45245\
        );

    \I__10584\ : SRMux
    port map (
            O => \N__45607\,
            I => \N__45245\
        );

    \I__10583\ : SRMux
    port map (
            O => \N__45606\,
            I => \N__45245\
        );

    \I__10582\ : SRMux
    port map (
            O => \N__45605\,
            I => \N__45245\
        );

    \I__10581\ : SRMux
    port map (
            O => \N__45604\,
            I => \N__45245\
        );

    \I__10580\ : SRMux
    port map (
            O => \N__45603\,
            I => \N__45245\
        );

    \I__10579\ : SRMux
    port map (
            O => \N__45602\,
            I => \N__45245\
        );

    \I__10578\ : SRMux
    port map (
            O => \N__45601\,
            I => \N__45245\
        );

    \I__10577\ : SRMux
    port map (
            O => \N__45600\,
            I => \N__45245\
        );

    \I__10576\ : SRMux
    port map (
            O => \N__45599\,
            I => \N__45245\
        );

    \I__10575\ : SRMux
    port map (
            O => \N__45598\,
            I => \N__45245\
        );

    \I__10574\ : SRMux
    port map (
            O => \N__45597\,
            I => \N__45245\
        );

    \I__10573\ : SRMux
    port map (
            O => \N__45596\,
            I => \N__45245\
        );

    \I__10572\ : SRMux
    port map (
            O => \N__45595\,
            I => \N__45245\
        );

    \I__10571\ : SRMux
    port map (
            O => \N__45594\,
            I => \N__45245\
        );

    \I__10570\ : SRMux
    port map (
            O => \N__45593\,
            I => \N__45245\
        );

    \I__10569\ : SRMux
    port map (
            O => \N__45592\,
            I => \N__45245\
        );

    \I__10568\ : SRMux
    port map (
            O => \N__45591\,
            I => \N__45245\
        );

    \I__10567\ : SRMux
    port map (
            O => \N__45590\,
            I => \N__45245\
        );

    \I__10566\ : SRMux
    port map (
            O => \N__45589\,
            I => \N__45245\
        );

    \I__10565\ : SRMux
    port map (
            O => \N__45588\,
            I => \N__45245\
        );

    \I__10564\ : SRMux
    port map (
            O => \N__45587\,
            I => \N__45245\
        );

    \I__10563\ : SRMux
    port map (
            O => \N__45586\,
            I => \N__45245\
        );

    \I__10562\ : SRMux
    port map (
            O => \N__45585\,
            I => \N__45245\
        );

    \I__10561\ : SRMux
    port map (
            O => \N__45584\,
            I => \N__45245\
        );

    \I__10560\ : SRMux
    port map (
            O => \N__45583\,
            I => \N__45245\
        );

    \I__10559\ : SRMux
    port map (
            O => \N__45582\,
            I => \N__45245\
        );

    \I__10558\ : SRMux
    port map (
            O => \N__45581\,
            I => \N__45245\
        );

    \I__10557\ : SRMux
    port map (
            O => \N__45580\,
            I => \N__45245\
        );

    \I__10556\ : SRMux
    port map (
            O => \N__45579\,
            I => \N__45245\
        );

    \I__10555\ : SRMux
    port map (
            O => \N__45578\,
            I => \N__45245\
        );

    \I__10554\ : SRMux
    port map (
            O => \N__45577\,
            I => \N__45245\
        );

    \I__10553\ : SRMux
    port map (
            O => \N__45576\,
            I => \N__45245\
        );

    \I__10552\ : SRMux
    port map (
            O => \N__45575\,
            I => \N__45245\
        );

    \I__10551\ : SRMux
    port map (
            O => \N__45574\,
            I => \N__45245\
        );

    \I__10550\ : SRMux
    port map (
            O => \N__45573\,
            I => \N__45245\
        );

    \I__10549\ : SRMux
    port map (
            O => \N__45572\,
            I => \N__45245\
        );

    \I__10548\ : SRMux
    port map (
            O => \N__45571\,
            I => \N__45245\
        );

    \I__10547\ : SRMux
    port map (
            O => \N__45570\,
            I => \N__45245\
        );

    \I__10546\ : SRMux
    port map (
            O => \N__45569\,
            I => \N__45245\
        );

    \I__10545\ : SRMux
    port map (
            O => \N__45568\,
            I => \N__45245\
        );

    \I__10544\ : SRMux
    port map (
            O => \N__45567\,
            I => \N__45245\
        );

    \I__10543\ : SRMux
    port map (
            O => \N__45566\,
            I => \N__45245\
        );

    \I__10542\ : SRMux
    port map (
            O => \N__45565\,
            I => \N__45245\
        );

    \I__10541\ : SRMux
    port map (
            O => \N__45564\,
            I => \N__45245\
        );

    \I__10540\ : SRMux
    port map (
            O => \N__45563\,
            I => \N__45245\
        );

    \I__10539\ : SRMux
    port map (
            O => \N__45562\,
            I => \N__45245\
        );

    \I__10538\ : SRMux
    port map (
            O => \N__45561\,
            I => \N__45245\
        );

    \I__10537\ : SRMux
    port map (
            O => \N__45560\,
            I => \N__45245\
        );

    \I__10536\ : SRMux
    port map (
            O => \N__45559\,
            I => \N__45245\
        );

    \I__10535\ : SRMux
    port map (
            O => \N__45558\,
            I => \N__45245\
        );

    \I__10534\ : SRMux
    port map (
            O => \N__45557\,
            I => \N__45245\
        );

    \I__10533\ : SRMux
    port map (
            O => \N__45556\,
            I => \N__45245\
        );

    \I__10532\ : SRMux
    port map (
            O => \N__45555\,
            I => \N__45245\
        );

    \I__10531\ : SRMux
    port map (
            O => \N__45554\,
            I => \N__45245\
        );

    \I__10530\ : SRMux
    port map (
            O => \N__45553\,
            I => \N__45245\
        );

    \I__10529\ : SRMux
    port map (
            O => \N__45552\,
            I => \N__45245\
        );

    \I__10528\ : SRMux
    port map (
            O => \N__45551\,
            I => \N__45245\
        );

    \I__10527\ : SRMux
    port map (
            O => \N__45550\,
            I => \N__45245\
        );

    \I__10526\ : SRMux
    port map (
            O => \N__45549\,
            I => \N__45245\
        );

    \I__10525\ : SRMux
    port map (
            O => \N__45548\,
            I => \N__45245\
        );

    \I__10524\ : SRMux
    port map (
            O => \N__45547\,
            I => \N__45245\
        );

    \I__10523\ : SRMux
    port map (
            O => \N__45546\,
            I => \N__45245\
        );

    \I__10522\ : SRMux
    port map (
            O => \N__45545\,
            I => \N__45245\
        );

    \I__10521\ : SRMux
    port map (
            O => \N__45544\,
            I => \N__45245\
        );

    \I__10520\ : SRMux
    port map (
            O => \N__45543\,
            I => \N__45245\
        );

    \I__10519\ : SRMux
    port map (
            O => \N__45542\,
            I => \N__45245\
        );

    \I__10518\ : SRMux
    port map (
            O => \N__45541\,
            I => \N__45245\
        );

    \I__10517\ : SRMux
    port map (
            O => \N__45540\,
            I => \N__45245\
        );

    \I__10516\ : SRMux
    port map (
            O => \N__45539\,
            I => \N__45245\
        );

    \I__10515\ : SRMux
    port map (
            O => \N__45538\,
            I => \N__45245\
        );

    \I__10514\ : SRMux
    port map (
            O => \N__45537\,
            I => \N__45245\
        );

    \I__10513\ : SRMux
    port map (
            O => \N__45536\,
            I => \N__45245\
        );

    \I__10512\ : SRMux
    port map (
            O => \N__45535\,
            I => \N__45245\
        );

    \I__10511\ : SRMux
    port map (
            O => \N__45534\,
            I => \N__45245\
        );

    \I__10510\ : SRMux
    port map (
            O => \N__45533\,
            I => \N__45245\
        );

    \I__10509\ : SRMux
    port map (
            O => \N__45532\,
            I => \N__45245\
        );

    \I__10508\ : SRMux
    port map (
            O => \N__45531\,
            I => \N__45245\
        );

    \I__10507\ : SRMux
    port map (
            O => \N__45530\,
            I => \N__45245\
        );

    \I__10506\ : SRMux
    port map (
            O => \N__45529\,
            I => \N__45245\
        );

    \I__10505\ : SRMux
    port map (
            O => \N__45528\,
            I => \N__45245\
        );

    \I__10504\ : SRMux
    port map (
            O => \N__45527\,
            I => \N__45245\
        );

    \I__10503\ : SRMux
    port map (
            O => \N__45526\,
            I => \N__45245\
        );

    \I__10502\ : Glb2LocalMux
    port map (
            O => \N__45523\,
            I => \N__45245\
        );

    \I__10501\ : Glb2LocalMux
    port map (
            O => \N__45520\,
            I => \N__45245\
        );

    \I__10500\ : SRMux
    port map (
            O => \N__45519\,
            I => \N__45245\
        );

    \I__10499\ : Glb2LocalMux
    port map (
            O => \N__45516\,
            I => \N__45245\
        );

    \I__10498\ : SRMux
    port map (
            O => \N__45515\,
            I => \N__45245\
        );

    \I__10497\ : SRMux
    port map (
            O => \N__45514\,
            I => \N__45245\
        );

    \I__10496\ : GlobalMux
    port map (
            O => \N__45245\,
            I => \N__45242\
        );

    \I__10495\ : gio2CtrlBuf
    port map (
            O => \N__45242\,
            I => red_c_g
        );

    \I__10494\ : CascadeMux
    port map (
            O => \N__45239\,
            I => \N__45235\
        );

    \I__10493\ : CascadeMux
    port map (
            O => \N__45238\,
            I => \N__45232\
        );

    \I__10492\ : InMux
    port map (
            O => \N__45235\,
            I => \N__45229\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45232\,
            I => \N__45225\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__45229\,
            I => \N__45221\
        );

    \I__10489\ : InMux
    port map (
            O => \N__45228\,
            I => \N__45218\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__45225\,
            I => \N__45215\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45224\,
            I => \N__45212\
        );

    \I__10486\ : Span4Mux_h
    port map (
            O => \N__45221\,
            I => \N__45209\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45218\,
            I => \N__45206\
        );

    \I__10484\ : Span4Mux_h
    port map (
            O => \N__45215\,
            I => \N__45201\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__45212\,
            I => \N__45201\
        );

    \I__10482\ : Span4Mux_v
    port map (
            O => \N__45209\,
            I => \N__45196\
        );

    \I__10481\ : Span4Mux_h
    port map (
            O => \N__45206\,
            I => \N__45196\
        );

    \I__10480\ : Odrv4
    port map (
            O => \N__45201\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10479\ : Odrv4
    port map (
            O => \N__45196\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10478\ : InMux
    port map (
            O => \N__45191\,
            I => \N__45187\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45190\,
            I => \N__45184\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__45187\,
            I => \N__45180\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__45184\,
            I => \N__45177\
        );

    \I__10474\ : InMux
    port map (
            O => \N__45183\,
            I => \N__45174\
        );

    \I__10473\ : Odrv12
    port map (
            O => \N__45180\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10472\ : Odrv4
    port map (
            O => \N__45177\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__45174\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10470\ : CascadeMux
    port map (
            O => \N__45167\,
            I => \N__45164\
        );

    \I__10469\ : InMux
    port map (
            O => \N__45164\,
            I => \N__45161\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__45161\,
            I => \N__45158\
        );

    \I__10467\ : Odrv12
    port map (
            O => \N__45158\,
            I => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\
        );

    \I__10466\ : CascadeMux
    port map (
            O => \N__45155\,
            I => \N__45151\
        );

    \I__10465\ : CascadeMux
    port map (
            O => \N__45154\,
            I => \N__45148\
        );

    \I__10464\ : InMux
    port map (
            O => \N__45151\,
            I => \N__45145\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45148\,
            I => \N__45142\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__45145\,
            I => \N__45138\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__45142\,
            I => \N__45135\
        );

    \I__10460\ : InMux
    port map (
            O => \N__45141\,
            I => \N__45132\
        );

    \I__10459\ : Span4Mux_h
    port map (
            O => \N__45138\,
            I => \N__45126\
        );

    \I__10458\ : Span4Mux_v
    port map (
            O => \N__45135\,
            I => \N__45126\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__45132\,
            I => \N__45123\
        );

    \I__10456\ : InMux
    port map (
            O => \N__45131\,
            I => \N__45120\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__45126\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10454\ : Odrv12
    port map (
            O => \N__45123\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__45120\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45113\,
            I => \N__45109\
        );

    \I__10451\ : InMux
    port map (
            O => \N__45112\,
            I => \N__45106\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__45109\,
            I => \N__45102\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__45106\,
            I => \N__45099\
        );

    \I__10448\ : InMux
    port map (
            O => \N__45105\,
            I => \N__45096\
        );

    \I__10447\ : Odrv12
    port map (
            O => \N__45102\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10446\ : Odrv4
    port map (
            O => \N__45099\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__45096\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45089\,
            I => \N__45086\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__45086\,
            I => \N__45083\
        );

    \I__10442\ : Odrv4
    port map (
            O => \N__45083\,
            I => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45080\,
            I => \N__45076\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45079\,
            I => \N__45072\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__45076\,
            I => \N__45069\
        );

    \I__10438\ : InMux
    port map (
            O => \N__45075\,
            I => \N__45066\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__45072\,
            I => \N__45061\
        );

    \I__10436\ : Span4Mux_v
    port map (
            O => \N__45069\,
            I => \N__45061\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__45066\,
            I => \N__45057\
        );

    \I__10434\ : Span4Mux_h
    port map (
            O => \N__45061\,
            I => \N__45054\
        );

    \I__10433\ : InMux
    port map (
            O => \N__45060\,
            I => \N__45051\
        );

    \I__10432\ : Span4Mux_h
    port map (
            O => \N__45057\,
            I => \N__45048\
        );

    \I__10431\ : Odrv4
    port map (
            O => \N__45054\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__45051\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10429\ : Odrv4
    port map (
            O => \N__45048\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10428\ : CascadeMux
    port map (
            O => \N__45041\,
            I => \N__45038\
        );

    \I__10427\ : InMux
    port map (
            O => \N__45038\,
            I => \N__45033\
        );

    \I__10426\ : InMux
    port map (
            O => \N__45037\,
            I => \N__45030\
        );

    \I__10425\ : InMux
    port map (
            O => \N__45036\,
            I => \N__45027\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__45033\,
            I => \N__45024\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__45030\,
            I => \N__45021\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__45027\,
            I => \N__45018\
        );

    \I__10421\ : Span4Mux_h
    port map (
            O => \N__45024\,
            I => \N__45015\
        );

    \I__10420\ : Span4Mux_h
    port map (
            O => \N__45021\,
            I => \N__45012\
        );

    \I__10419\ : Odrv4
    port map (
            O => \N__45018\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10418\ : Odrv4
    port map (
            O => \N__45015\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10417\ : Odrv4
    port map (
            O => \N__45012\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45005\,
            I => \N__45002\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__45002\,
            I => \N__44999\
        );

    \I__10414\ : Odrv4
    port map (
            O => \N__44999\,
            I => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\
        );

    \I__10413\ : CascadeMux
    port map (
            O => \N__44996\,
            I => \N__44993\
        );

    \I__10412\ : InMux
    port map (
            O => \N__44993\,
            I => \N__44990\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__44990\,
            I => \N__44987\
        );

    \I__10410\ : Span4Mux_h
    port map (
            O => \N__44987\,
            I => \N__44983\
        );

    \I__10409\ : InMux
    port map (
            O => \N__44986\,
            I => \N__44980\
        );

    \I__10408\ : Span4Mux_v
    port map (
            O => \N__44983\,
            I => \N__44975\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__44980\,
            I => \N__44972\
        );

    \I__10406\ : InMux
    port map (
            O => \N__44979\,
            I => \N__44969\
        );

    \I__10405\ : InMux
    port map (
            O => \N__44978\,
            I => \N__44966\
        );

    \I__10404\ : Odrv4
    port map (
            O => \N__44975\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__10403\ : Odrv12
    port map (
            O => \N__44972\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__44969\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__44966\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__10400\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44954\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__44954\,
            I => \N__44949\
        );

    \I__10398\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44946\
        );

    \I__10397\ : CascadeMux
    port map (
            O => \N__44952\,
            I => \N__44943\
        );

    \I__10396\ : Span4Mux_v
    port map (
            O => \N__44949\,
            I => \N__44938\
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__44946\,
            I => \N__44938\
        );

    \I__10394\ : InMux
    port map (
            O => \N__44943\,
            I => \N__44935\
        );

    \I__10393\ : Span4Mux_h
    port map (
            O => \N__44938\,
            I => \N__44932\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__44935\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__10391\ : Odrv4
    port map (
            O => \N__44932\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__10390\ : InMux
    port map (
            O => \N__44927\,
            I => \N__44924\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__44924\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__10388\ : CascadeMux
    port map (
            O => \N__44921\,
            I => \N__44918\
        );

    \I__10387\ : InMux
    port map (
            O => \N__44918\,
            I => \N__44912\
        );

    \I__10386\ : InMux
    port map (
            O => \N__44917\,
            I => \N__44905\
        );

    \I__10385\ : InMux
    port map (
            O => \N__44916\,
            I => \N__44905\
        );

    \I__10384\ : InMux
    port map (
            O => \N__44915\,
            I => \N__44905\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__44912\,
            I => \N__44902\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__44905\,
            I => \N__44899\
        );

    \I__10381\ : Span4Mux_v
    port map (
            O => \N__44902\,
            I => \N__44896\
        );

    \I__10380\ : Span4Mux_h
    port map (
            O => \N__44899\,
            I => \N__44893\
        );

    \I__10379\ : Span4Mux_v
    port map (
            O => \N__44896\,
            I => \N__44888\
        );

    \I__10378\ : Span4Mux_v
    port map (
            O => \N__44893\,
            I => \N__44888\
        );

    \I__10377\ : Odrv4
    port map (
            O => \N__44888\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__10376\ : InMux
    port map (
            O => \N__44885\,
            I => \N__44882\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__44882\,
            I => \N__44879\
        );

    \I__10374\ : Span4Mux_h
    port map (
            O => \N__44879\,
            I => \N__44874\
        );

    \I__10373\ : InMux
    port map (
            O => \N__44878\,
            I => \N__44869\
        );

    \I__10372\ : InMux
    port map (
            O => \N__44877\,
            I => \N__44869\
        );

    \I__10371\ : Odrv4
    port map (
            O => \N__44874\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__44869\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__10369\ : InMux
    port map (
            O => \N__44864\,
            I => \N__44861\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__44861\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__10367\ : CascadeMux
    port map (
            O => \N__44858\,
            I => \N__44854\
        );

    \I__10366\ : CascadeMux
    port map (
            O => \N__44857\,
            I => \N__44851\
        );

    \I__10365\ : InMux
    port map (
            O => \N__44854\,
            I => \N__44848\
        );

    \I__10364\ : InMux
    port map (
            O => \N__44851\,
            I => \N__44845\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__44848\,
            I => \N__44842\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__44845\,
            I => \N__44837\
        );

    \I__10361\ : Span4Mux_v
    port map (
            O => \N__44842\,
            I => \N__44834\
        );

    \I__10360\ : InMux
    port map (
            O => \N__44841\,
            I => \N__44831\
        );

    \I__10359\ : InMux
    port map (
            O => \N__44840\,
            I => \N__44828\
        );

    \I__10358\ : Odrv12
    port map (
            O => \N__44837\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10357\ : Odrv4
    port map (
            O => \N__44834\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__44831\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__44828\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10354\ : InMux
    port map (
            O => \N__44819\,
            I => \N__44815\
        );

    \I__10353\ : InMux
    port map (
            O => \N__44818\,
            I => \N__44812\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__44815\,
            I => \N__44808\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__44812\,
            I => \N__44805\
        );

    \I__10350\ : InMux
    port map (
            O => \N__44811\,
            I => \N__44802\
        );

    \I__10349\ : Span4Mux_h
    port map (
            O => \N__44808\,
            I => \N__44797\
        );

    \I__10348\ : Span4Mux_v
    port map (
            O => \N__44805\,
            I => \N__44797\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__44802\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__10346\ : Odrv4
    port map (
            O => \N__44797\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__10345\ : CascadeMux
    port map (
            O => \N__44792\,
            I => \N__44789\
        );

    \I__10344\ : InMux
    port map (
            O => \N__44789\,
            I => \N__44786\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__44786\,
            I => \N__44783\
        );

    \I__10342\ : Odrv4
    port map (
            O => \N__44783\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__10341\ : CascadeMux
    port map (
            O => \N__44780\,
            I => \N__44777\
        );

    \I__10340\ : InMux
    port map (
            O => \N__44777\,
            I => \N__44772\
        );

    \I__10339\ : CascadeMux
    port map (
            O => \N__44776\,
            I => \N__44769\
        );

    \I__10338\ : InMux
    port map (
            O => \N__44775\,
            I => \N__44766\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__44772\,
            I => \N__44763\
        );

    \I__10336\ : InMux
    port map (
            O => \N__44769\,
            I => \N__44760\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__44766\,
            I => \N__44757\
        );

    \I__10334\ : Span12Mux_v
    port map (
            O => \N__44763\,
            I => \N__44753\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__44760\,
            I => \N__44750\
        );

    \I__10332\ : Span4Mux_v
    port map (
            O => \N__44757\,
            I => \N__44747\
        );

    \I__10331\ : InMux
    port map (
            O => \N__44756\,
            I => \N__44744\
        );

    \I__10330\ : Odrv12
    port map (
            O => \N__44753\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10329\ : Odrv12
    port map (
            O => \N__44750\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10328\ : Odrv4
    port map (
            O => \N__44747\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__44744\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10326\ : InMux
    port map (
            O => \N__44735\,
            I => \N__44730\
        );

    \I__10325\ : InMux
    port map (
            O => \N__44734\,
            I => \N__44727\
        );

    \I__10324\ : InMux
    port map (
            O => \N__44733\,
            I => \N__44724\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__44730\,
            I => \N__44719\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__44727\,
            I => \N__44719\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__44724\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10320\ : Odrv12
    port map (
            O => \N__44719\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10319\ : InMux
    port map (
            O => \N__44714\,
            I => \N__44711\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__44711\,
            I => \N__44708\
        );

    \I__10317\ : Odrv4
    port map (
            O => \N__44708\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__10316\ : CascadeMux
    port map (
            O => \N__44705\,
            I => \N__44702\
        );

    \I__10315\ : InMux
    port map (
            O => \N__44702\,
            I => \N__44699\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__44699\,
            I => \N__44694\
        );

    \I__10313\ : InMux
    port map (
            O => \N__44698\,
            I => \N__44691\
        );

    \I__10312\ : InMux
    port map (
            O => \N__44697\,
            I => \N__44688\
        );

    \I__10311\ : Odrv12
    port map (
            O => \N__44694\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__44691\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__44688\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__10308\ : InMux
    port map (
            O => \N__44681\,
            I => \N__44676\
        );

    \I__10307\ : InMux
    port map (
            O => \N__44680\,
            I => \N__44673\
        );

    \I__10306\ : InMux
    port map (
            O => \N__44679\,
            I => \N__44670\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__44676\,
            I => \N__44667\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__44673\,
            I => \N__44664\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__44670\,
            I => \N__44660\
        );

    \I__10302\ : Span4Mux_v
    port map (
            O => \N__44667\,
            I => \N__44655\
        );

    \I__10301\ : Span4Mux_v
    port map (
            O => \N__44664\,
            I => \N__44655\
        );

    \I__10300\ : InMux
    port map (
            O => \N__44663\,
            I => \N__44652\
        );

    \I__10299\ : Odrv4
    port map (
            O => \N__44660\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10298\ : Odrv4
    port map (
            O => \N__44655\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__44652\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10296\ : CascadeMux
    port map (
            O => \N__44645\,
            I => \N__44642\
        );

    \I__10295\ : InMux
    port map (
            O => \N__44642\,
            I => \N__44639\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__44639\,
            I => \N__44636\
        );

    \I__10293\ : Span4Mux_h
    port map (
            O => \N__44636\,
            I => \N__44633\
        );

    \I__10292\ : Odrv4
    port map (
            O => \N__44633\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__10291\ : InMux
    port map (
            O => \N__44630\,
            I => \N__44627\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__44627\,
            I => \N__44624\
        );

    \I__10289\ : Span4Mux_h
    port map (
            O => \N__44624\,
            I => \N__44621\
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__44621\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__10287\ : InMux
    port map (
            O => \N__44618\,
            I => \bfn_18_17_0_\
        );

    \I__10286\ : InMux
    port map (
            O => \N__44615\,
            I => \N__44612\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__44612\,
            I => \N__44609\
        );

    \I__10284\ : Span4Mux_h
    port map (
            O => \N__44609\,
            I => \N__44606\
        );

    \I__10283\ : Odrv4
    port map (
            O => \N__44606\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__10282\ : InMux
    port map (
            O => \N__44603\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__10281\ : CascadeMux
    port map (
            O => \N__44600\,
            I => \N__44597\
        );

    \I__10280\ : InMux
    port map (
            O => \N__44597\,
            I => \N__44594\
        );

    \I__10279\ : LocalMux
    port map (
            O => \N__44594\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__10278\ : InMux
    port map (
            O => \N__44591\,
            I => \N__44588\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__44588\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__10276\ : InMux
    port map (
            O => \N__44585\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__10275\ : InMux
    port map (
            O => \N__44582\,
            I => \N__44579\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__44579\,
            I => \N__44576\
        );

    \I__10273\ : Span4Mux_h
    port map (
            O => \N__44576\,
            I => \N__44573\
        );

    \I__10272\ : Odrv4
    port map (
            O => \N__44573\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__10271\ : InMux
    port map (
            O => \N__44570\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__10270\ : CascadeMux
    port map (
            O => \N__44567\,
            I => \N__44564\
        );

    \I__10269\ : InMux
    port map (
            O => \N__44564\,
            I => \N__44561\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__44561\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__10267\ : InMux
    port map (
            O => \N__44558\,
            I => \N__44555\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__44555\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__10265\ : InMux
    port map (
            O => \N__44552\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__10264\ : InMux
    port map (
            O => \N__44549\,
            I => \N__44546\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__44546\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__10262\ : InMux
    port map (
            O => \N__44543\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__10261\ : CascadeMux
    port map (
            O => \N__44540\,
            I => \N__44536\
        );

    \I__10260\ : CascadeMux
    port map (
            O => \N__44539\,
            I => \N__44533\
        );

    \I__10259\ : InMux
    port map (
            O => \N__44536\,
            I => \N__44530\
        );

    \I__10258\ : InMux
    port map (
            O => \N__44533\,
            I => \N__44527\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__44530\,
            I => \N__44524\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__44527\,
            I => \N__44519\
        );

    \I__10255\ : Span4Mux_h
    port map (
            O => \N__44524\,
            I => \N__44519\
        );

    \I__10254\ : Odrv4
    port map (
            O => \N__44519\,
            I => \current_shift_inst.un4_control_input_0_31\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44516\,
            I => \N__44513\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__44513\,
            I => \N__44510\
        );

    \I__10251\ : Span4Mux_h
    port map (
            O => \N__44510\,
            I => \N__44507\
        );

    \I__10250\ : Odrv4
    port map (
            O => \N__44507\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__10249\ : InMux
    port map (
            O => \N__44504\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__10248\ : InMux
    port map (
            O => \N__44501\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__10247\ : CascadeMux
    port map (
            O => \N__44498\,
            I => \N__44495\
        );

    \I__10246\ : InMux
    port map (
            O => \N__44495\,
            I => \N__44492\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__44492\,
            I => \N__44489\
        );

    \I__10244\ : Odrv4
    port map (
            O => \N__44489\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44486\,
            I => \N__44483\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__44483\,
            I => \N__44480\
        );

    \I__10241\ : Odrv4
    port map (
            O => \N__44480\,
            I => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\
        );

    \I__10240\ : CascadeMux
    port map (
            O => \N__44477\,
            I => \N__44474\
        );

    \I__10239\ : InMux
    port map (
            O => \N__44474\,
            I => \N__44471\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__44471\,
            I => \N__44468\
        );

    \I__10237\ : Span4Mux_h
    port map (
            O => \N__44468\,
            I => \N__44465\
        );

    \I__10236\ : Span4Mux_h
    port map (
            O => \N__44465\,
            I => \N__44462\
        );

    \I__10235\ : Odrv4
    port map (
            O => \N__44462\,
            I => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\
        );

    \I__10234\ : InMux
    port map (
            O => \N__44459\,
            I => \N__44456\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__44456\,
            I => \N__44453\
        );

    \I__10232\ : Span4Mux_h
    port map (
            O => \N__44453\,
            I => \N__44450\
        );

    \I__10231\ : Odrv4
    port map (
            O => \N__44450\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__10230\ : InMux
    port map (
            O => \N__44447\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__10229\ : InMux
    port map (
            O => \N__44444\,
            I => \N__44441\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__44441\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__10227\ : InMux
    port map (
            O => \N__44438\,
            I => \N__44435\
        );

    \I__10226\ : LocalMux
    port map (
            O => \N__44435\,
            I => \N__44432\
        );

    \I__10225\ : Odrv4
    port map (
            O => \N__44432\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__10224\ : InMux
    port map (
            O => \N__44429\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__10223\ : CascadeMux
    port map (
            O => \N__44426\,
            I => \N__44423\
        );

    \I__10222\ : InMux
    port map (
            O => \N__44423\,
            I => \N__44420\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__44420\,
            I => \N__44417\
        );

    \I__10220\ : Span4Mux_h
    port map (
            O => \N__44417\,
            I => \N__44414\
        );

    \I__10219\ : Odrv4
    port map (
            O => \N__44414\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__10218\ : InMux
    port map (
            O => \N__44411\,
            I => \N__44408\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__44408\,
            I => \N__44405\
        );

    \I__10216\ : Odrv12
    port map (
            O => \N__44405\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__10215\ : InMux
    port map (
            O => \N__44402\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__10214\ : InMux
    port map (
            O => \N__44399\,
            I => \N__44396\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__44396\,
            I => \N__44393\
        );

    \I__10212\ : Span4Mux_h
    port map (
            O => \N__44393\,
            I => \N__44390\
        );

    \I__10211\ : Odrv4
    port map (
            O => \N__44390\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__10210\ : InMux
    port map (
            O => \N__44387\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__10209\ : InMux
    port map (
            O => \N__44384\,
            I => \N__44381\
        );

    \I__10208\ : LocalMux
    port map (
            O => \N__44381\,
            I => \N__44378\
        );

    \I__10207\ : Odrv4
    port map (
            O => \N__44378\,
            I => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\
        );

    \I__10206\ : CascadeMux
    port map (
            O => \N__44375\,
            I => \N__44372\
        );

    \I__10205\ : InMux
    port map (
            O => \N__44372\,
            I => \N__44369\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__44369\,
            I => \N__44366\
        );

    \I__10203\ : Span4Mux_h
    port map (
            O => \N__44366\,
            I => \N__44363\
        );

    \I__10202\ : Odrv4
    port map (
            O => \N__44363\,
            I => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\
        );

    \I__10201\ : InMux
    port map (
            O => \N__44360\,
            I => \N__44357\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__44357\,
            I => \N__44354\
        );

    \I__10199\ : Span4Mux_h
    port map (
            O => \N__44354\,
            I => \N__44351\
        );

    \I__10198\ : Odrv4
    port map (
            O => \N__44351\,
            I => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\
        );

    \I__10197\ : CascadeMux
    port map (
            O => \N__44348\,
            I => \N__44345\
        );

    \I__10196\ : InMux
    port map (
            O => \N__44345\,
            I => \N__44342\
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__44342\,
            I => \N__44339\
        );

    \I__10194\ : Odrv12
    port map (
            O => \N__44339\,
            I => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\
        );

    \I__10193\ : CascadeMux
    port map (
            O => \N__44336\,
            I => \N__44333\
        );

    \I__10192\ : InMux
    port map (
            O => \N__44333\,
            I => \N__44330\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__44330\,
            I => \N__44327\
        );

    \I__10190\ : Span4Mux_h
    port map (
            O => \N__44327\,
            I => \N__44324\
        );

    \I__10189\ : Odrv4
    port map (
            O => \N__44324\,
            I => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\
        );

    \I__10188\ : CascadeMux
    port map (
            O => \N__44321\,
            I => \N__44318\
        );

    \I__10187\ : InMux
    port map (
            O => \N__44318\,
            I => \N__44315\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__44315\,
            I => \N__44312\
        );

    \I__10185\ : Span4Mux_v
    port map (
            O => \N__44312\,
            I => \N__44309\
        );

    \I__10184\ : Odrv4
    port map (
            O => \N__44309\,
            I => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\
        );

    \I__10183\ : InMux
    port map (
            O => \N__44306\,
            I => \N__44303\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__44303\,
            I => \N__44300\
        );

    \I__10181\ : Span4Mux_h
    port map (
            O => \N__44300\,
            I => \N__44297\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__44297\,
            I => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\
        );

    \I__10179\ : CEMux
    port map (
            O => \N__44294\,
            I => \N__44286\
        );

    \I__10178\ : CEMux
    port map (
            O => \N__44293\,
            I => \N__44283\
        );

    \I__10177\ : CEMux
    port map (
            O => \N__44292\,
            I => \N__44280\
        );

    \I__10176\ : CEMux
    port map (
            O => \N__44291\,
            I => \N__44277\
        );

    \I__10175\ : CEMux
    port map (
            O => \N__44290\,
            I => \N__44274\
        );

    \I__10174\ : CEMux
    port map (
            O => \N__44289\,
            I => \N__44253\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__44286\,
            I => \N__44250\
        );

    \I__10172\ : LocalMux
    port map (
            O => \N__44283\,
            I => \N__44247\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__44280\,
            I => \N__44244\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__44277\,
            I => \N__44238\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__44274\,
            I => \N__44238\
        );

    \I__10168\ : InMux
    port map (
            O => \N__44273\,
            I => \N__44231\
        );

    \I__10167\ : InMux
    port map (
            O => \N__44272\,
            I => \N__44231\
        );

    \I__10166\ : InMux
    port map (
            O => \N__44271\,
            I => \N__44231\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44270\,
            I => \N__44228\
        );

    \I__10164\ : InMux
    port map (
            O => \N__44269\,
            I => \N__44223\
        );

    \I__10163\ : InMux
    port map (
            O => \N__44268\,
            I => \N__44223\
        );

    \I__10162\ : InMux
    port map (
            O => \N__44267\,
            I => \N__44214\
        );

    \I__10161\ : InMux
    port map (
            O => \N__44266\,
            I => \N__44214\
        );

    \I__10160\ : InMux
    port map (
            O => \N__44265\,
            I => \N__44214\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44264\,
            I => \N__44214\
        );

    \I__10158\ : InMux
    port map (
            O => \N__44263\,
            I => \N__44205\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44262\,
            I => \N__44205\
        );

    \I__10156\ : InMux
    port map (
            O => \N__44261\,
            I => \N__44205\
        );

    \I__10155\ : InMux
    port map (
            O => \N__44260\,
            I => \N__44205\
        );

    \I__10154\ : InMux
    port map (
            O => \N__44259\,
            I => \N__44196\
        );

    \I__10153\ : InMux
    port map (
            O => \N__44258\,
            I => \N__44196\
        );

    \I__10152\ : InMux
    port map (
            O => \N__44257\,
            I => \N__44196\
        );

    \I__10151\ : InMux
    port map (
            O => \N__44256\,
            I => \N__44196\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__44253\,
            I => \N__44193\
        );

    \I__10149\ : Span4Mux_v
    port map (
            O => \N__44250\,
            I => \N__44188\
        );

    \I__10148\ : Span4Mux_h
    port map (
            O => \N__44247\,
            I => \N__44188\
        );

    \I__10147\ : Span4Mux_v
    port map (
            O => \N__44244\,
            I => \N__44185\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44243\,
            I => \N__44182\
        );

    \I__10145\ : Span4Mux_v
    port map (
            O => \N__44238\,
            I => \N__44179\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__44231\,
            I => \N__44176\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__44228\,
            I => \N__44165\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__44223\,
            I => \N__44165\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__44214\,
            I => \N__44165\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__44205\,
            I => \N__44165\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__44196\,
            I => \N__44165\
        );

    \I__10138\ : Span4Mux_v
    port map (
            O => \N__44193\,
            I => \N__44160\
        );

    \I__10137\ : Span4Mux_v
    port map (
            O => \N__44188\,
            I => \N__44160\
        );

    \I__10136\ : Span4Mux_h
    port map (
            O => \N__44185\,
            I => \N__44155\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__44182\,
            I => \N__44155\
        );

    \I__10134\ : Span4Mux_v
    port map (
            O => \N__44179\,
            I => \N__44148\
        );

    \I__10133\ : Span4Mux_v
    port map (
            O => \N__44176\,
            I => \N__44148\
        );

    \I__10132\ : Span4Mux_v
    port map (
            O => \N__44165\,
            I => \N__44148\
        );

    \I__10131\ : Odrv4
    port map (
            O => \N__44160\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__10130\ : Odrv4
    port map (
            O => \N__44155\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__10129\ : Odrv4
    port map (
            O => \N__44148\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44141\,
            I => \N__44134\
        );

    \I__10127\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44134\
        );

    \I__10126\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44131\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__44134\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__10124\ : LocalMux
    port map (
            O => \N__44131\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__10123\ : CascadeMux
    port map (
            O => \N__44126\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\
        );

    \I__10122\ : CascadeMux
    port map (
            O => \N__44123\,
            I => \N__44118\
        );

    \I__10121\ : InMux
    port map (
            O => \N__44122\,
            I => \N__44115\
        );

    \I__10120\ : InMux
    port map (
            O => \N__44121\,
            I => \N__44112\
        );

    \I__10119\ : InMux
    port map (
            O => \N__44118\,
            I => \N__44109\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__44115\,
            I => \N__44106\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__44112\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__44109\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10115\ : Odrv4
    port map (
            O => \N__44106\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10114\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44096\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__44096\,
            I => \N__44092\
        );

    \I__10112\ : CascadeMux
    port map (
            O => \N__44095\,
            I => \N__44089\
        );

    \I__10111\ : Span4Mux_h
    port map (
            O => \N__44092\,
            I => \N__44086\
        );

    \I__10110\ : InMux
    port map (
            O => \N__44089\,
            I => \N__44083\
        );

    \I__10109\ : Odrv4
    port map (
            O => \N__44086\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__44083\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__10107\ : InMux
    port map (
            O => \N__44078\,
            I => \N__44074\
        );

    \I__10106\ : CascadeMux
    port map (
            O => \N__44077\,
            I => \N__44071\
        );

    \I__10105\ : LocalMux
    port map (
            O => \N__44074\,
            I => \N__44068\
        );

    \I__10104\ : InMux
    port map (
            O => \N__44071\,
            I => \N__44065\
        );

    \I__10103\ : Span4Mux_v
    port map (
            O => \N__44068\,
            I => \N__44062\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44065\,
            I => \N__44059\
        );

    \I__10101\ : Odrv4
    port map (
            O => \N__44062\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__10100\ : Odrv12
    port map (
            O => \N__44059\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__10099\ : CascadeMux
    port map (
            O => \N__44054\,
            I => \N__44050\
        );

    \I__10098\ : InMux
    port map (
            O => \N__44053\,
            I => \N__44045\
        );

    \I__10097\ : InMux
    port map (
            O => \N__44050\,
            I => \N__44045\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__44045\,
            I => \N__44041\
        );

    \I__10095\ : InMux
    port map (
            O => \N__44044\,
            I => \N__44037\
        );

    \I__10094\ : Span4Mux_v
    port map (
            O => \N__44041\,
            I => \N__44034\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44040\,
            I => \N__44031\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__44037\,
            I => \N__44028\
        );

    \I__10091\ : Odrv4
    port map (
            O => \N__44034\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__44031\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10089\ : Odrv12
    port map (
            O => \N__44028\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10088\ : CascadeMux
    port map (
            O => \N__44021\,
            I => \N__44018\
        );

    \I__10087\ : InMux
    port map (
            O => \N__44018\,
            I => \N__44015\
        );

    \I__10086\ : LocalMux
    port map (
            O => \N__44015\,
            I => \N__44012\
        );

    \I__10085\ : Span4Mux_h
    port map (
            O => \N__44012\,
            I => \N__44009\
        );

    \I__10084\ : Span4Mux_h
    port map (
            O => \N__44009\,
            I => \N__44006\
        );

    \I__10083\ : Odrv4
    port map (
            O => \N__44006\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__10082\ : CascadeMux
    port map (
            O => \N__44003\,
            I => \N__44000\
        );

    \I__10081\ : InMux
    port map (
            O => \N__44000\,
            I => \N__43997\
        );

    \I__10080\ : LocalMux
    port map (
            O => \N__43997\,
            I => \N__43994\
        );

    \I__10079\ : Span4Mux_h
    port map (
            O => \N__43994\,
            I => \N__43991\
        );

    \I__10078\ : Odrv4
    port map (
            O => \N__43991\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__10077\ : InMux
    port map (
            O => \N__43988\,
            I => \N__43985\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__43985\,
            I => \N__43982\
        );

    \I__10075\ : Span4Mux_v
    port map (
            O => \N__43982\,
            I => \N__43979\
        );

    \I__10074\ : Odrv4
    port map (
            O => \N__43979\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__10073\ : CascadeMux
    port map (
            O => \N__43976\,
            I => \N__43973\
        );

    \I__10072\ : InMux
    port map (
            O => \N__43973\,
            I => \N__43970\
        );

    \I__10071\ : LocalMux
    port map (
            O => \N__43970\,
            I => \N__43967\
        );

    \I__10070\ : Span4Mux_h
    port map (
            O => \N__43967\,
            I => \N__43964\
        );

    \I__10069\ : Odrv4
    port map (
            O => \N__43964\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__10068\ : InMux
    port map (
            O => \N__43961\,
            I => \N__43958\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__43958\,
            I => \N__43955\
        );

    \I__10066\ : Span4Mux_h
    port map (
            O => \N__43955\,
            I => \N__43952\
        );

    \I__10065\ : Span4Mux_h
    port map (
            O => \N__43952\,
            I => \N__43949\
        );

    \I__10064\ : Odrv4
    port map (
            O => \N__43949\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__10063\ : CascadeMux
    port map (
            O => \N__43946\,
            I => \N__43943\
        );

    \I__10062\ : InMux
    port map (
            O => \N__43943\,
            I => \N__43940\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__43940\,
            I => \N__43937\
        );

    \I__10060\ : Odrv12
    port map (
            O => \N__43937\,
            I => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\
        );

    \I__10059\ : InMux
    port map (
            O => \N__43934\,
            I => \N__43930\
        );

    \I__10058\ : InMux
    port map (
            O => \N__43933\,
            I => \N__43927\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__43930\,
            I => \N__43922\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__43927\,
            I => \N__43919\
        );

    \I__10055\ : InMux
    port map (
            O => \N__43926\,
            I => \N__43916\
        );

    \I__10054\ : InMux
    port map (
            O => \N__43925\,
            I => \N__43913\
        );

    \I__10053\ : Span12Mux_s7_h
    port map (
            O => \N__43922\,
            I => \N__43908\
        );

    \I__10052\ : Span12Mux_s9_v
    port map (
            O => \N__43919\,
            I => \N__43908\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__43916\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__43913\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__10049\ : Odrv12
    port map (
            O => \N__43908\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__10048\ : InMux
    port map (
            O => \N__43901\,
            I => \N__43898\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__43898\,
            I => \N__43892\
        );

    \I__10046\ : InMux
    port map (
            O => \N__43897\,
            I => \N__43889\
        );

    \I__10045\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43884\
        );

    \I__10044\ : InMux
    port map (
            O => \N__43895\,
            I => \N__43884\
        );

    \I__10043\ : Span4Mux_h
    port map (
            O => \N__43892\,
            I => \N__43881\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__43889\,
            I => \N__43878\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__43884\,
            I => \N__43874\
        );

    \I__10040\ : Span4Mux_v
    port map (
            O => \N__43881\,
            I => \N__43869\
        );

    \I__10039\ : Span4Mux_h
    port map (
            O => \N__43878\,
            I => \N__43869\
        );

    \I__10038\ : InMux
    port map (
            O => \N__43877\,
            I => \N__43866\
        );

    \I__10037\ : Span4Mux_h
    port map (
            O => \N__43874\,
            I => \N__43863\
        );

    \I__10036\ : Span4Mux_h
    port map (
            O => \N__43869\,
            I => \N__43860\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__43866\,
            I => \N__43855\
        );

    \I__10034\ : Span4Mux_h
    port map (
            O => \N__43863\,
            I => \N__43855\
        );

    \I__10033\ : Odrv4
    port map (
            O => \N__43860\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__10032\ : Odrv4
    port map (
            O => \N__43855\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__10031\ : CascadeMux
    port map (
            O => \N__43850\,
            I => \N__43847\
        );

    \I__10030\ : InMux
    port map (
            O => \N__43847\,
            I => \N__43842\
        );

    \I__10029\ : InMux
    port map (
            O => \N__43846\,
            I => \N__43839\
        );

    \I__10028\ : InMux
    port map (
            O => \N__43845\,
            I => \N__43836\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__43842\,
            I => \N__43832\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__43839\,
            I => \N__43829\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__43836\,
            I => \N__43826\
        );

    \I__10024\ : CascadeMux
    port map (
            O => \N__43835\,
            I => \N__43822\
        );

    \I__10023\ : Span4Mux_v
    port map (
            O => \N__43832\,
            I => \N__43817\
        );

    \I__10022\ : Span4Mux_v
    port map (
            O => \N__43829\,
            I => \N__43817\
        );

    \I__10021\ : Span4Mux_h
    port map (
            O => \N__43826\,
            I => \N__43814\
        );

    \I__10020\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43811\
        );

    \I__10019\ : InMux
    port map (
            O => \N__43822\,
            I => \N__43808\
        );

    \I__10018\ : Span4Mux_h
    port map (
            O => \N__43817\,
            I => \N__43805\
        );

    \I__10017\ : Span4Mux_h
    port map (
            O => \N__43814\,
            I => \N__43800\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__43811\,
            I => \N__43800\
        );

    \I__10015\ : LocalMux
    port map (
            O => \N__43808\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__10014\ : Odrv4
    port map (
            O => \N__43805\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__10013\ : Odrv4
    port map (
            O => \N__43800\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__10012\ : InMux
    port map (
            O => \N__43793\,
            I => \N__43789\
        );

    \I__10011\ : InMux
    port map (
            O => \N__43792\,
            I => \N__43786\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__43789\,
            I => \N__43783\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__43786\,
            I => \N__43777\
        );

    \I__10008\ : Span4Mux_h
    port map (
            O => \N__43783\,
            I => \N__43777\
        );

    \I__10007\ : InMux
    port map (
            O => \N__43782\,
            I => \N__43774\
        );

    \I__10006\ : Span4Mux_h
    port map (
            O => \N__43777\,
            I => \N__43769\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__43774\,
            I => \N__43769\
        );

    \I__10004\ : Span4Mux_v
    port map (
            O => \N__43769\,
            I => \N__43766\
        );

    \I__10003\ : Odrv4
    port map (
            O => \N__43766\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO\
        );

    \I__10002\ : InMux
    port map (
            O => \N__43763\,
            I => \N__43759\
        );

    \I__10001\ : InMux
    port map (
            O => \N__43762\,
            I => \N__43756\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__43759\,
            I => \N__43753\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__43756\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__9998\ : Odrv4
    port map (
            O => \N__43753\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__9997\ : InMux
    port map (
            O => \N__43748\,
            I => \N__43745\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__43745\,
            I => \N__43742\
        );

    \I__9995\ : Span4Mux_h
    port map (
            O => \N__43742\,
            I => \N__43737\
        );

    \I__9994\ : InMux
    port map (
            O => \N__43741\,
            I => \N__43734\
        );

    \I__9993\ : InMux
    port map (
            O => \N__43740\,
            I => \N__43731\
        );

    \I__9992\ : Span4Mux_h
    port map (
            O => \N__43737\,
            I => \N__43728\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__43734\,
            I => \N__43725\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__43731\,
            I => \N__43722\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__43728\,
            I => \N__43719\
        );

    \I__9988\ : Span4Mux_v
    port map (
            O => \N__43725\,
            I => \N__43716\
        );

    \I__9987\ : Span4Mux_v
    port map (
            O => \N__43722\,
            I => \N__43713\
        );

    \I__9986\ : Sp12to4
    port map (
            O => \N__43719\,
            I => \N__43710\
        );

    \I__9985\ : Span4Mux_h
    port map (
            O => \N__43716\,
            I => \N__43707\
        );

    \I__9984\ : Odrv4
    port map (
            O => \N__43713\,
            I => \il_min_comp2_D2\
        );

    \I__9983\ : Odrv12
    port map (
            O => \N__43710\,
            I => \il_min_comp2_D2\
        );

    \I__9982\ : Odrv4
    port map (
            O => \N__43707\,
            I => \il_min_comp2_D2\
        );

    \I__9981\ : InMux
    port map (
            O => \N__43700\,
            I => \N__43697\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__43697\,
            I => \phase_controller_inst2.start_timer_tr_0_sqmuxa\
        );

    \I__9979\ : InMux
    port map (
            O => \N__43694\,
            I => \N__43691\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__43691\,
            I => \N__43688\
        );

    \I__9977\ : Span4Mux_h
    port map (
            O => \N__43688\,
            I => \N__43685\
        );

    \I__9976\ : Span4Mux_h
    port map (
            O => \N__43685\,
            I => \N__43682\
        );

    \I__9975\ : Odrv4
    port map (
            O => \N__43682\,
            I => \phase_controller_inst2.time_passed_RNI9M3O\
        );

    \I__9974\ : CascadeMux
    port map (
            O => \N__43679\,
            I => \N__43674\
        );

    \I__9973\ : CascadeMux
    port map (
            O => \N__43678\,
            I => \N__43671\
        );

    \I__9972\ : InMux
    port map (
            O => \N__43677\,
            I => \N__43668\
        );

    \I__9971\ : InMux
    port map (
            O => \N__43674\,
            I => \N__43665\
        );

    \I__9970\ : InMux
    port map (
            O => \N__43671\,
            I => \N__43660\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__43668\,
            I => \N__43657\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__43665\,
            I => \N__43654\
        );

    \I__9967\ : InMux
    port map (
            O => \N__43664\,
            I => \N__43651\
        );

    \I__9966\ : InMux
    port map (
            O => \N__43663\,
            I => \N__43647\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__43660\,
            I => \N__43644\
        );

    \I__9964\ : Span4Mux_v
    port map (
            O => \N__43657\,
            I => \N__43641\
        );

    \I__9963\ : Span4Mux_h
    port map (
            O => \N__43654\,
            I => \N__43636\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__43651\,
            I => \N__43636\
        );

    \I__9961\ : InMux
    port map (
            O => \N__43650\,
            I => \N__43633\
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__43647\,
            I => \N__43628\
        );

    \I__9959\ : Span4Mux_h
    port map (
            O => \N__43644\,
            I => \N__43628\
        );

    \I__9958\ : Span4Mux_v
    port map (
            O => \N__43641\,
            I => \N__43623\
        );

    \I__9957\ : Span4Mux_h
    port map (
            O => \N__43636\,
            I => \N__43623\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__43633\,
            I => phase_controller_inst1_state_4
        );

    \I__9955\ : Odrv4
    port map (
            O => \N__43628\,
            I => phase_controller_inst1_state_4
        );

    \I__9954\ : Odrv4
    port map (
            O => \N__43623\,
            I => phase_controller_inst1_state_4
        );

    \I__9953\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43613\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__43613\,
            I => \N__43609\
        );

    \I__9951\ : InMux
    port map (
            O => \N__43612\,
            I => \N__43605\
        );

    \I__9950\ : Span4Mux_h
    port map (
            O => \N__43609\,
            I => \N__43602\
        );

    \I__9949\ : InMux
    port map (
            O => \N__43608\,
            I => \N__43599\
        );

    \I__9948\ : LocalMux
    port map (
            O => \N__43605\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO\
        );

    \I__9947\ : Odrv4
    port map (
            O => \N__43602\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__43599\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO\
        );

    \I__9945\ : CascadeMux
    port map (
            O => \N__43592\,
            I => \N__43589\
        );

    \I__9944\ : InMux
    port map (
            O => \N__43589\,
            I => \N__43586\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__43586\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLHZ0Z1\
        );

    \I__9942\ : CascadeMux
    port map (
            O => \N__43583\,
            I => \N__43580\
        );

    \I__9941\ : InMux
    port map (
            O => \N__43580\,
            I => \N__43577\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__43577\,
            I => \N__43574\
        );

    \I__9939\ : Span4Mux_h
    port map (
            O => \N__43574\,
            I => \N__43569\
        );

    \I__9938\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43566\
        );

    \I__9937\ : CascadeMux
    port map (
            O => \N__43572\,
            I => \N__43562\
        );

    \I__9936\ : Span4Mux_h
    port map (
            O => \N__43569\,
            I => \N__43558\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__43566\,
            I => \N__43555\
        );

    \I__9934\ : InMux
    port map (
            O => \N__43565\,
            I => \N__43552\
        );

    \I__9933\ : InMux
    port map (
            O => \N__43562\,
            I => \N__43547\
        );

    \I__9932\ : InMux
    port map (
            O => \N__43561\,
            I => \N__43547\
        );

    \I__9931\ : Odrv4
    port map (
            O => \N__43558\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__9930\ : Odrv4
    port map (
            O => \N__43555\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__43552\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__43547\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__9927\ : InMux
    port map (
            O => \N__43538\,
            I => \N__43532\
        );

    \I__9926\ : InMux
    port map (
            O => \N__43537\,
            I => \N__43532\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__43532\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__9924\ : InMux
    port map (
            O => \N__43529\,
            I => \N__43526\
        );

    \I__9923\ : LocalMux
    port map (
            O => \N__43526\,
            I => \N__43520\
        );

    \I__9922\ : InMux
    port map (
            O => \N__43525\,
            I => \N__43513\
        );

    \I__9921\ : InMux
    port map (
            O => \N__43524\,
            I => \N__43513\
        );

    \I__9920\ : InMux
    port map (
            O => \N__43523\,
            I => \N__43513\
        );

    \I__9919\ : Odrv12
    port map (
            O => \N__43520\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__43513\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__9917\ : InMux
    port map (
            O => \N__43508\,
            I => \N__43505\
        );

    \I__9916\ : LocalMux
    port map (
            O => \N__43505\,
            I => \N__43502\
        );

    \I__9915\ : Span4Mux_h
    port map (
            O => \N__43502\,
            I => \N__43499\
        );

    \I__9914\ : Span4Mux_h
    port map (
            O => \N__43499\,
            I => \N__43493\
        );

    \I__9913\ : InMux
    port map (
            O => \N__43498\,
            I => \N__43488\
        );

    \I__9912\ : InMux
    port map (
            O => \N__43497\,
            I => \N__43488\
        );

    \I__9911\ : InMux
    port map (
            O => \N__43496\,
            I => \N__43485\
        );

    \I__9910\ : Odrv4
    port map (
            O => \N__43493\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__43488\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__43485\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__9907\ : CascadeMux
    port map (
            O => \N__43478\,
            I => \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\
        );

    \I__9906\ : InMux
    port map (
            O => \N__43475\,
            I => \N__43471\
        );

    \I__9905\ : InMux
    port map (
            O => \N__43474\,
            I => \N__43468\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__43471\,
            I => \elapsed_time_ns_1_RNI0GIF91_0_26\
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__43468\,
            I => \elapsed_time_ns_1_RNI0GIF91_0_26\
        );

    \I__9902\ : InMux
    port map (
            O => \N__43463\,
            I => \N__43460\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__43460\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15\
        );

    \I__9900\ : InMux
    port map (
            O => \N__43457\,
            I => \N__43454\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__43454\,
            I => \N__43450\
        );

    \I__9898\ : InMux
    port map (
            O => \N__43453\,
            I => \N__43447\
        );

    \I__9897\ : Span4Mux_h
    port map (
            O => \N__43450\,
            I => \N__43442\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__43447\,
            I => \N__43442\
        );

    \I__9895\ : Odrv4
    port map (
            O => \N__43442\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__9894\ : InMux
    port map (
            O => \N__43439\,
            I => \N__43433\
        );

    \I__9893\ : InMux
    port map (
            O => \N__43438\,
            I => \N__43433\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__43433\,
            I => \elapsed_time_ns_1_RNI2IIF91_0_28\
        );

    \I__9891\ : InMux
    port map (
            O => \N__43430\,
            I => \N__43423\
        );

    \I__9890\ : InMux
    port map (
            O => \N__43429\,
            I => \N__43420\
        );

    \I__9889\ : InMux
    port map (
            O => \N__43428\,
            I => \N__43417\
        );

    \I__9888\ : InMux
    port map (
            O => \N__43427\,
            I => \N__43414\
        );

    \I__9887\ : InMux
    port map (
            O => \N__43426\,
            I => \N__43411\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__43423\,
            I => \N__43408\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__43420\,
            I => \N__43405\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__43417\,
            I => \N__43398\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__43414\,
            I => \N__43398\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__43411\,
            I => \N__43398\
        );

    \I__9881\ : Span4Mux_v
    port map (
            O => \N__43408\,
            I => \N__43393\
        );

    \I__9880\ : Span4Mux_v
    port map (
            O => \N__43405\,
            I => \N__43393\
        );

    \I__9879\ : Span4Mux_h
    port map (
            O => \N__43398\,
            I => \N__43390\
        );

    \I__9878\ : Odrv4
    port map (
            O => \N__43393\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__9877\ : Odrv4
    port map (
            O => \N__43390\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__9876\ : CascadeMux
    port map (
            O => \N__43385\,
            I => \N__43382\
        );

    \I__9875\ : InMux
    port map (
            O => \N__43382\,
            I => \N__43379\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__43379\,
            I => \N__43374\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43378\,
            I => \N__43369\
        );

    \I__9872\ : InMux
    port map (
            O => \N__43377\,
            I => \N__43369\
        );

    \I__9871\ : Span4Mux_h
    port map (
            O => \N__43374\,
            I => \N__43366\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__43369\,
            I => \delay_measurement_inst.delay_tr_timer.N_378\
        );

    \I__9869\ : Odrv4
    port map (
            O => \N__43366\,
            I => \delay_measurement_inst.delay_tr_timer.N_378\
        );

    \I__9868\ : InMux
    port map (
            O => \N__43361\,
            I => \N__43358\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__43358\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0\
        );

    \I__9866\ : InMux
    port map (
            O => \N__43355\,
            I => \N__43352\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__43352\,
            I => \N__43348\
        );

    \I__9864\ : InMux
    port map (
            O => \N__43351\,
            I => \N__43345\
        );

    \I__9863\ : Odrv4
    port map (
            O => \N__43348\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__43345\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__9861\ : CascadeMux
    port map (
            O => \N__43340\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\
        );

    \I__9860\ : InMux
    port map (
            O => \N__43337\,
            I => \N__43333\
        );

    \I__9859\ : InMux
    port map (
            O => \N__43336\,
            I => \N__43330\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__43333\,
            I => \N__43324\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__43330\,
            I => \N__43324\
        );

    \I__9856\ : InMux
    port map (
            O => \N__43329\,
            I => \N__43320\
        );

    \I__9855\ : Span4Mux_v
    port map (
            O => \N__43324\,
            I => \N__43317\
        );

    \I__9854\ : InMux
    port map (
            O => \N__43323\,
            I => \N__43314\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__43320\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__9852\ : Odrv4
    port map (
            O => \N__43317\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__43314\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__9850\ : InMux
    port map (
            O => \N__43307\,
            I => \N__43303\
        );

    \I__9849\ : CascadeMux
    port map (
            O => \N__43306\,
            I => \N__43300\
        );

    \I__9848\ : LocalMux
    port map (
            O => \N__43303\,
            I => \N__43297\
        );

    \I__9847\ : InMux
    port map (
            O => \N__43300\,
            I => \N__43294\
        );

    \I__9846\ : Span4Mux_h
    port map (
            O => \N__43297\,
            I => \N__43289\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__43294\,
            I => \N__43289\
        );

    \I__9844\ : Odrv4
    port map (
            O => \N__43289\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__9843\ : CascadeMux
    port map (
            O => \N__43286\,
            I => \N__43283\
        );

    \I__9842\ : InMux
    port map (
            O => \N__43283\,
            I => \N__43280\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__43280\,
            I => \N__43276\
        );

    \I__9840\ : InMux
    port map (
            O => \N__43279\,
            I => \N__43273\
        );

    \I__9839\ : Odrv4
    port map (
            O => \N__43276\,
            I => \elapsed_time_ns_1_RNI1HIF91_0_27\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__43273\,
            I => \elapsed_time_ns_1_RNI1HIF91_0_27\
        );

    \I__9837\ : InMux
    port map (
            O => \N__43268\,
            I => \N__43264\
        );

    \I__9836\ : CascadeMux
    port map (
            O => \N__43267\,
            I => \N__43261\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__43264\,
            I => \N__43258\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43261\,
            I => \N__43255\
        );

    \I__9833\ : Span4Mux_v
    port map (
            O => \N__43258\,
            I => \N__43252\
        );

    \I__9832\ : LocalMux
    port map (
            O => \N__43255\,
            I => \N__43249\
        );

    \I__9831\ : Odrv4
    port map (
            O => \N__43252\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9830\ : Odrv4
    port map (
            O => \N__43249\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9829\ : CascadeMux
    port map (
            O => \N__43244\,
            I => \N__43241\
        );

    \I__9828\ : InMux
    port map (
            O => \N__43241\,
            I => \N__43237\
        );

    \I__9827\ : InMux
    port map (
            O => \N__43240\,
            I => \N__43234\
        );

    \I__9826\ : LocalMux
    port map (
            O => \N__43237\,
            I => \elapsed_time_ns_1_RNISBIF91_0_22\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__43234\,
            I => \elapsed_time_ns_1_RNISBIF91_0_22\
        );

    \I__9824\ : InMux
    port map (
            O => \N__43229\,
            I => \N__43225\
        );

    \I__9823\ : InMux
    port map (
            O => \N__43228\,
            I => \N__43222\
        );

    \I__9822\ : LocalMux
    port map (
            O => \N__43225\,
            I => \N__43219\
        );

    \I__9821\ : LocalMux
    port map (
            O => \N__43222\,
            I => \N__43216\
        );

    \I__9820\ : Span4Mux_v
    port map (
            O => \N__43219\,
            I => \N__43213\
        );

    \I__9819\ : Span4Mux_h
    port map (
            O => \N__43216\,
            I => \N__43210\
        );

    \I__9818\ : Odrv4
    port map (
            O => \N__43213\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9817\ : Odrv4
    port map (
            O => \N__43210\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43205\,
            I => \N__43201\
        );

    \I__9815\ : InMux
    port map (
            O => \N__43204\,
            I => \N__43198\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__43201\,
            I => \elapsed_time_ns_1_RNIQ9IF91_0_20\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__43198\,
            I => \elapsed_time_ns_1_RNIQ9IF91_0_20\
        );

    \I__9812\ : InMux
    port map (
            O => \N__43193\,
            I => \N__43190\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__43190\,
            I => \N__43186\
        );

    \I__9810\ : InMux
    port map (
            O => \N__43189\,
            I => \N__43183\
        );

    \I__9809\ : Span4Mux_v
    port map (
            O => \N__43186\,
            I => \N__43180\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__43183\,
            I => \N__43177\
        );

    \I__9807\ : Odrv4
    port map (
            O => \N__43180\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9806\ : Odrv4
    port map (
            O => \N__43177\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9805\ : CascadeMux
    port map (
            O => \N__43172\,
            I => \N__43164\
        );

    \I__9804\ : CascadeMux
    port map (
            O => \N__43171\,
            I => \N__43161\
        );

    \I__9803\ : CascadeMux
    port map (
            O => \N__43170\,
            I => \N__43158\
        );

    \I__9802\ : CascadeMux
    port map (
            O => \N__43169\,
            I => \N__43153\
        );

    \I__9801\ : InMux
    port map (
            O => \N__43168\,
            I => \N__43149\
        );

    \I__9800\ : InMux
    port map (
            O => \N__43167\,
            I => \N__43142\
        );

    \I__9799\ : InMux
    port map (
            O => \N__43164\,
            I => \N__43134\
        );

    \I__9798\ : InMux
    port map (
            O => \N__43161\,
            I => \N__43127\
        );

    \I__9797\ : InMux
    port map (
            O => \N__43158\,
            I => \N__43127\
        );

    \I__9796\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43127\
        );

    \I__9795\ : InMux
    port map (
            O => \N__43156\,
            I => \N__43122\
        );

    \I__9794\ : InMux
    port map (
            O => \N__43153\,
            I => \N__43122\
        );

    \I__9793\ : InMux
    port map (
            O => \N__43152\,
            I => \N__43118\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__43149\,
            I => \N__43115\
        );

    \I__9791\ : InMux
    port map (
            O => \N__43148\,
            I => \N__43108\
        );

    \I__9790\ : InMux
    port map (
            O => \N__43147\,
            I => \N__43108\
        );

    \I__9789\ : InMux
    port map (
            O => \N__43146\,
            I => \N__43108\
        );

    \I__9788\ : CascadeMux
    port map (
            O => \N__43145\,
            I => \N__43104\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__43142\,
            I => \N__43096\
        );

    \I__9786\ : InMux
    port map (
            O => \N__43141\,
            I => \N__43093\
        );

    \I__9785\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43090\
        );

    \I__9784\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43085\
        );

    \I__9783\ : InMux
    port map (
            O => \N__43138\,
            I => \N__43085\
        );

    \I__9782\ : InMux
    port map (
            O => \N__43137\,
            I => \N__43082\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__43134\,
            I => \N__43079\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__43127\,
            I => \N__43074\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__43122\,
            I => \N__43074\
        );

    \I__9778\ : CascadeMux
    port map (
            O => \N__43121\,
            I => \N__43066\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__43118\,
            I => \N__43059\
        );

    \I__9776\ : Span4Mux_v
    port map (
            O => \N__43115\,
            I => \N__43059\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__43108\,
            I => \N__43059\
        );

    \I__9774\ : InMux
    port map (
            O => \N__43107\,
            I => \N__43052\
        );

    \I__9773\ : InMux
    port map (
            O => \N__43104\,
            I => \N__43052\
        );

    \I__9772\ : InMux
    port map (
            O => \N__43103\,
            I => \N__43052\
        );

    \I__9771\ : InMux
    port map (
            O => \N__43102\,
            I => \N__43049\
        );

    \I__9770\ : InMux
    port map (
            O => \N__43101\,
            I => \N__43042\
        );

    \I__9769\ : InMux
    port map (
            O => \N__43100\,
            I => \N__43042\
        );

    \I__9768\ : InMux
    port map (
            O => \N__43099\,
            I => \N__43042\
        );

    \I__9767\ : Span4Mux_h
    port map (
            O => \N__43096\,
            I => \N__43031\
        );

    \I__9766\ : LocalMux
    port map (
            O => \N__43093\,
            I => \N__43031\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__43090\,
            I => \N__43031\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__43085\,
            I => \N__43031\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__43082\,
            I => \N__43031\
        );

    \I__9762\ : Span4Mux_h
    port map (
            O => \N__43079\,
            I => \N__43026\
        );

    \I__9761\ : Span4Mux_v
    port map (
            O => \N__43074\,
            I => \N__43026\
        );

    \I__9760\ : InMux
    port map (
            O => \N__43073\,
            I => \N__43013\
        );

    \I__9759\ : InMux
    port map (
            O => \N__43072\,
            I => \N__43013\
        );

    \I__9758\ : InMux
    port map (
            O => \N__43071\,
            I => \N__43013\
        );

    \I__9757\ : InMux
    port map (
            O => \N__43070\,
            I => \N__43013\
        );

    \I__9756\ : InMux
    port map (
            O => \N__43069\,
            I => \N__43013\
        );

    \I__9755\ : InMux
    port map (
            O => \N__43066\,
            I => \N__43013\
        );

    \I__9754\ : Span4Mux_h
    port map (
            O => \N__43059\,
            I => \N__43008\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__43052\,
            I => \N__43008\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__43049\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__43042\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9750\ : Odrv4
    port map (
            O => \N__43031\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9749\ : Odrv4
    port map (
            O => \N__43026\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__43013\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9747\ : Odrv4
    port map (
            O => \N__43008\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9746\ : CascadeMux
    port map (
            O => \N__42995\,
            I => \N__42987\
        );

    \I__9745\ : CascadeMux
    port map (
            O => \N__42994\,
            I => \N__42984\
        );

    \I__9744\ : InMux
    port map (
            O => \N__42993\,
            I => \N__42979\
        );

    \I__9743\ : CascadeMux
    port map (
            O => \N__42992\,
            I => \N__42976\
        );

    \I__9742\ : CascadeMux
    port map (
            O => \N__42991\,
            I => \N__42972\
        );

    \I__9741\ : InMux
    port map (
            O => \N__42990\,
            I => \N__42968\
        );

    \I__9740\ : InMux
    port map (
            O => \N__42987\,
            I => \N__42963\
        );

    \I__9739\ : InMux
    port map (
            O => \N__42984\,
            I => \N__42963\
        );

    \I__9738\ : CascadeMux
    port map (
            O => \N__42983\,
            I => \N__42959\
        );

    \I__9737\ : CascadeMux
    port map (
            O => \N__42982\,
            I => \N__42953\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__42979\,
            I => \N__42947\
        );

    \I__9735\ : InMux
    port map (
            O => \N__42976\,
            I => \N__42944\
        );

    \I__9734\ : CascadeMux
    port map (
            O => \N__42975\,
            I => \N__42937\
        );

    \I__9733\ : InMux
    port map (
            O => \N__42972\,
            I => \N__42934\
        );

    \I__9732\ : InMux
    port map (
            O => \N__42971\,
            I => \N__42931\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__42968\,
            I => \N__42926\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__42963\,
            I => \N__42926\
        );

    \I__9729\ : InMux
    port map (
            O => \N__42962\,
            I => \N__42923\
        );

    \I__9728\ : InMux
    port map (
            O => \N__42959\,
            I => \N__42916\
        );

    \I__9727\ : InMux
    port map (
            O => \N__42958\,
            I => \N__42916\
        );

    \I__9726\ : InMux
    port map (
            O => \N__42957\,
            I => \N__42916\
        );

    \I__9725\ : InMux
    port map (
            O => \N__42956\,
            I => \N__42913\
        );

    \I__9724\ : InMux
    port map (
            O => \N__42953\,
            I => \N__42908\
        );

    \I__9723\ : InMux
    port map (
            O => \N__42952\,
            I => \N__42908\
        );

    \I__9722\ : InMux
    port map (
            O => \N__42951\,
            I => \N__42903\
        );

    \I__9721\ : InMux
    port map (
            O => \N__42950\,
            I => \N__42903\
        );

    \I__9720\ : Span4Mux_h
    port map (
            O => \N__42947\,
            I => \N__42898\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__42944\,
            I => \N__42898\
        );

    \I__9718\ : InMux
    port map (
            O => \N__42943\,
            I => \N__42889\
        );

    \I__9717\ : InMux
    port map (
            O => \N__42942\,
            I => \N__42889\
        );

    \I__9716\ : InMux
    port map (
            O => \N__42941\,
            I => \N__42889\
        );

    \I__9715\ : InMux
    port map (
            O => \N__42940\,
            I => \N__42889\
        );

    \I__9714\ : InMux
    port map (
            O => \N__42937\,
            I => \N__42886\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__42934\,
            I => \N__42881\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__42931\,
            I => \N__42881\
        );

    \I__9711\ : Span4Mux_v
    port map (
            O => \N__42926\,
            I => \N__42878\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__42923\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__42916\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__42913\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__9707\ : LocalMux
    port map (
            O => \N__42908\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__9706\ : LocalMux
    port map (
            O => \N__42903\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__9705\ : Odrv4
    port map (
            O => \N__42898\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__42889\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__42886\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__9702\ : Odrv12
    port map (
            O => \N__42881\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__9701\ : Odrv4
    port map (
            O => \N__42878\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__9700\ : CascadeMux
    port map (
            O => \N__42857\,
            I => \N__42854\
        );

    \I__9699\ : InMux
    port map (
            O => \N__42854\,
            I => \N__42850\
        );

    \I__9698\ : InMux
    port map (
            O => \N__42853\,
            I => \N__42847\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__42850\,
            I => \elapsed_time_ns_1_RNIRBJF91_0_30\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__42847\,
            I => \elapsed_time_ns_1_RNIRBJF91_0_30\
        );

    \I__9695\ : CascadeMux
    port map (
            O => \N__42842\,
            I => \N__42839\
        );

    \I__9694\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42835\
        );

    \I__9693\ : InMux
    port map (
            O => \N__42838\,
            I => \N__42832\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__42835\,
            I => \N__42827\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__42832\,
            I => \N__42827\
        );

    \I__9690\ : Odrv4
    port map (
            O => \N__42827\,
            I => \delay_measurement_inst.delay_tr_timer.N_367\
        );

    \I__9689\ : InMux
    port map (
            O => \N__42824\,
            I => \N__42820\
        );

    \I__9688\ : InMux
    port map (
            O => \N__42823\,
            I => \N__42817\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__42820\,
            I => \N__42814\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__42817\,
            I => \N__42811\
        );

    \I__9685\ : Span4Mux_v
    port map (
            O => \N__42814\,
            I => \N__42807\
        );

    \I__9684\ : Span4Mux_h
    port map (
            O => \N__42811\,
            I => \N__42804\
        );

    \I__9683\ : InMux
    port map (
            O => \N__42810\,
            I => \N__42801\
        );

    \I__9682\ : Odrv4
    port map (
            O => \N__42807\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__9681\ : Odrv4
    port map (
            O => \N__42804\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__42801\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__9679\ : CascadeMux
    port map (
            O => \N__42794\,
            I => \N__42791\
        );

    \I__9678\ : InMux
    port map (
            O => \N__42791\,
            I => \N__42786\
        );

    \I__9677\ : CascadeMux
    port map (
            O => \N__42790\,
            I => \N__42782\
        );

    \I__9676\ : CascadeMux
    port map (
            O => \N__42789\,
            I => \N__42779\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__42786\,
            I => \N__42776\
        );

    \I__9674\ : InMux
    port map (
            O => \N__42785\,
            I => \N__42771\
        );

    \I__9673\ : InMux
    port map (
            O => \N__42782\,
            I => \N__42771\
        );

    \I__9672\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42768\
        );

    \I__9671\ : Span4Mux_v
    port map (
            O => \N__42776\,
            I => \N__42765\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__42771\,
            I => \N__42762\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__42768\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__9668\ : Odrv4
    port map (
            O => \N__42765\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__9667\ : Odrv4
    port map (
            O => \N__42762\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__9666\ : InMux
    port map (
            O => \N__42755\,
            I => \N__42752\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__42752\,
            I => \delay_measurement_inst.delay_tr_timer.N_349\
        );

    \I__9664\ : CascadeMux
    port map (
            O => \N__42749\,
            I => \delay_measurement_inst.delay_tr_timer.N_363_cascade_\
        );

    \I__9663\ : CascadeMux
    port map (
            O => \N__42746\,
            I => \N__42742\
        );

    \I__9662\ : CascadeMux
    port map (
            O => \N__42745\,
            I => \N__42738\
        );

    \I__9661\ : InMux
    port map (
            O => \N__42742\,
            I => \N__42730\
        );

    \I__9660\ : InMux
    port map (
            O => \N__42741\,
            I => \N__42727\
        );

    \I__9659\ : InMux
    port map (
            O => \N__42738\,
            I => \N__42724\
        );

    \I__9658\ : InMux
    port map (
            O => \N__42737\,
            I => \N__42721\
        );

    \I__9657\ : InMux
    port map (
            O => \N__42736\,
            I => \N__42716\
        );

    \I__9656\ : InMux
    port map (
            O => \N__42735\,
            I => \N__42716\
        );

    \I__9655\ : InMux
    port map (
            O => \N__42734\,
            I => \N__42713\
        );

    \I__9654\ : InMux
    port map (
            O => \N__42733\,
            I => \N__42710\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__42730\,
            I => \N__42699\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__42727\,
            I => \N__42699\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__42724\,
            I => \N__42699\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__42721\,
            I => \N__42699\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__42716\,
            I => \N__42699\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__42713\,
            I => \N__42696\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__42710\,
            I => \N__42690\
        );

    \I__9646\ : Span4Mux_v
    port map (
            O => \N__42699\,
            I => \N__42690\
        );

    \I__9645\ : Span4Mux_v
    port map (
            O => \N__42696\,
            I => \N__42687\
        );

    \I__9644\ : InMux
    port map (
            O => \N__42695\,
            I => \N__42684\
        );

    \I__9643\ : Span4Mux_h
    port map (
            O => \N__42690\,
            I => \N__42681\
        );

    \I__9642\ : Odrv4
    port map (
            O => \N__42687\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__42684\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__9640\ : Odrv4
    port map (
            O => \N__42681\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__9639\ : InMux
    port map (
            O => \N__42674\,
            I => \N__42671\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__42671\,
            I => \N__42667\
        );

    \I__9637\ : InMux
    port map (
            O => \N__42670\,
            I => \N__42664\
        );

    \I__9636\ : Odrv4
    port map (
            O => \N__42667\,
            I => \delay_measurement_inst.delay_tr_timer.N_380\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__42664\,
            I => \delay_measurement_inst.delay_tr_timer.N_380\
        );

    \I__9634\ : CascadeMux
    port map (
            O => \N__42659\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_\
        );

    \I__9633\ : InMux
    port map (
            O => \N__42656\,
            I => \N__42653\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__42653\,
            I => \N__42650\
        );

    \I__9631\ : Odrv4
    port map (
            O => \N__42650\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6\
        );

    \I__9630\ : CascadeMux
    port map (
            O => \N__42647\,
            I => \N__42644\
        );

    \I__9629\ : InMux
    port map (
            O => \N__42644\,
            I => \N__42640\
        );

    \I__9628\ : InMux
    port map (
            O => \N__42643\,
            I => \N__42637\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__42640\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__42637\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\
        );

    \I__9625\ : InMux
    port map (
            O => \N__42632\,
            I => \N__42627\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42631\,
            I => \N__42622\
        );

    \I__9623\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42622\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__42627\,
            I => \N__42617\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__42622\,
            I => \N__42617\
        );

    \I__9620\ : Odrv4
    port map (
            O => \N__42617\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\
        );

    \I__9619\ : InMux
    port map (
            O => \N__42614\,
            I => \N__42609\
        );

    \I__9618\ : InMux
    port map (
            O => \N__42613\,
            I => \N__42604\
        );

    \I__9617\ : InMux
    port map (
            O => \N__42612\,
            I => \N__42604\
        );

    \I__9616\ : LocalMux
    port map (
            O => \N__42609\,
            I => \delay_measurement_inst.delay_tr_timer.N_365\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__42604\,
            I => \delay_measurement_inst.delay_tr_timer.N_365\
        );

    \I__9614\ : CascadeMux
    port map (
            O => \N__42599\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8_cascade_\
        );

    \I__9613\ : CascadeMux
    port map (
            O => \N__42596\,
            I => \N__42592\
        );

    \I__9612\ : InMux
    port map (
            O => \N__42595\,
            I => \N__42589\
        );

    \I__9611\ : InMux
    port map (
            O => \N__42592\,
            I => \N__42586\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__42589\,
            I => \delay_measurement_inst.delay_tr_timer.N_345\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__42586\,
            I => \delay_measurement_inst.delay_tr_timer.N_345\
        );

    \I__9608\ : InMux
    port map (
            O => \N__42581\,
            I => \N__42575\
        );

    \I__9607\ : InMux
    port map (
            O => \N__42580\,
            I => \N__42575\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__42575\,
            I => \delay_measurement_inst.delay_tr_timer.N_359_1\
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__42572\,
            I => \N__42568\
        );

    \I__9604\ : CascadeMux
    port map (
            O => \N__42571\,
            I => \N__42565\
        );

    \I__9603\ : InMux
    port map (
            O => \N__42568\,
            I => \N__42560\
        );

    \I__9602\ : InMux
    port map (
            O => \N__42565\,
            I => \N__42560\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__42560\,
            I => \N__42557\
        );

    \I__9600\ : Span4Mux_h
    port map (
            O => \N__42557\,
            I => \N__42554\
        );

    \I__9599\ : Odrv4
    port map (
            O => \N__42554\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9598\ : InMux
    port map (
            O => \N__42551\,
            I => \N__42548\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__42548\,
            I => \N__42545\
        );

    \I__9596\ : Span4Mux_v
    port map (
            O => \N__42545\,
            I => \N__42541\
        );

    \I__9595\ : InMux
    port map (
            O => \N__42544\,
            I => \N__42538\
        );

    \I__9594\ : Odrv4
    port map (
            O => \N__42541\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__42538\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__9592\ : CascadeMux
    port map (
            O => \N__42533\,
            I => \N__42530\
        );

    \I__9591\ : InMux
    port map (
            O => \N__42530\,
            I => \N__42526\
        );

    \I__9590\ : InMux
    port map (
            O => \N__42529\,
            I => \N__42523\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__42526\,
            I => \elapsed_time_ns_1_RNIUDIF91_0_24\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__42523\,
            I => \elapsed_time_ns_1_RNIUDIF91_0_24\
        );

    \I__9587\ : InMux
    port map (
            O => \N__42518\,
            I => \N__42514\
        );

    \I__9586\ : InMux
    port map (
            O => \N__42517\,
            I => \N__42511\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__42514\,
            I => \N__42508\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__42511\,
            I => \N__42505\
        );

    \I__9583\ : Span4Mux_h
    port map (
            O => \N__42508\,
            I => \N__42502\
        );

    \I__9582\ : Span4Mux_h
    port map (
            O => \N__42505\,
            I => \N__42499\
        );

    \I__9581\ : Odrv4
    port map (
            O => \N__42502\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__9580\ : Odrv4
    port map (
            O => \N__42499\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__9579\ : InMux
    port map (
            O => \N__42494\,
            I => \N__42491\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__42491\,
            I => \elapsed_time_ns_1_RNIVEIF91_0_25\
        );

    \I__9577\ : InMux
    port map (
            O => \N__42488\,
            I => \N__42483\
        );

    \I__9576\ : InMux
    port map (
            O => \N__42487\,
            I => \N__42480\
        );

    \I__9575\ : InMux
    port map (
            O => \N__42486\,
            I => \N__42477\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__42483\,
            I => \N__42474\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__42480\,
            I => \N__42471\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__42477\,
            I => \N__42468\
        );

    \I__9571\ : Span4Mux_h
    port map (
            O => \N__42474\,
            I => \N__42464\
        );

    \I__9570\ : Sp12to4
    port map (
            O => \N__42471\,
            I => \N__42461\
        );

    \I__9569\ : Span4Mux_h
    port map (
            O => \N__42468\,
            I => \N__42458\
        );

    \I__9568\ : InMux
    port map (
            O => \N__42467\,
            I => \N__42455\
        );

    \I__9567\ : Odrv4
    port map (
            O => \N__42464\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9566\ : Odrv12
    port map (
            O => \N__42461\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9565\ : Odrv4
    port map (
            O => \N__42458\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__42455\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9563\ : CascadeMux
    port map (
            O => \N__42446\,
            I => \N__42442\
        );

    \I__9562\ : CascadeMux
    port map (
            O => \N__42445\,
            I => \N__42438\
        );

    \I__9561\ : InMux
    port map (
            O => \N__42442\,
            I => \N__42435\
        );

    \I__9560\ : InMux
    port map (
            O => \N__42441\,
            I => \N__42432\
        );

    \I__9559\ : InMux
    port map (
            O => \N__42438\,
            I => \N__42429\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__42435\,
            I => \N__42426\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__42432\,
            I => \N__42423\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__42429\,
            I => \N__42420\
        );

    \I__9555\ : Span4Mux_h
    port map (
            O => \N__42426\,
            I => \N__42415\
        );

    \I__9554\ : Span4Mux_v
    port map (
            O => \N__42423\,
            I => \N__42415\
        );

    \I__9553\ : Odrv4
    port map (
            O => \N__42420\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9552\ : Odrv4
    port map (
            O => \N__42415\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9551\ : CascadeMux
    port map (
            O => \N__42410\,
            I => \N__42407\
        );

    \I__9550\ : InMux
    port map (
            O => \N__42407\,
            I => \N__42404\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__42404\,
            I => \N__42401\
        );

    \I__9548\ : Span4Mux_v
    port map (
            O => \N__42401\,
            I => \N__42398\
        );

    \I__9547\ : Odrv4
    port map (
            O => \N__42398\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42395\,
            I => \N__42391\
        );

    \I__9545\ : InMux
    port map (
            O => \N__42394\,
            I => \N__42388\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__42391\,
            I => \N__42383\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__42388\,
            I => \N__42380\
        );

    \I__9542\ : InMux
    port map (
            O => \N__42387\,
            I => \N__42377\
        );

    \I__9541\ : InMux
    port map (
            O => \N__42386\,
            I => \N__42374\
        );

    \I__9540\ : Span4Mux_v
    port map (
            O => \N__42383\,
            I => \N__42371\
        );

    \I__9539\ : Span4Mux_v
    port map (
            O => \N__42380\,
            I => \N__42368\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__42377\,
            I => \N__42365\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__42374\,
            I => \N__42362\
        );

    \I__9536\ : Odrv4
    port map (
            O => \N__42371\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9535\ : Odrv4
    port map (
            O => \N__42368\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9534\ : Odrv4
    port map (
            O => \N__42365\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9533\ : Odrv4
    port map (
            O => \N__42362\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9532\ : InMux
    port map (
            O => \N__42353\,
            I => \N__42350\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__42350\,
            I => \N__42347\
        );

    \I__9530\ : Span4Mux_h
    port map (
            O => \N__42347\,
            I => \N__42344\
        );

    \I__9529\ : Odrv4
    port map (
            O => \N__42344\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__9528\ : CascadeMux
    port map (
            O => \N__42341\,
            I => \N__42337\
        );

    \I__9527\ : CascadeMux
    port map (
            O => \N__42340\,
            I => \N__42334\
        );

    \I__9526\ : InMux
    port map (
            O => \N__42337\,
            I => \N__42331\
        );

    \I__9525\ : InMux
    port map (
            O => \N__42334\,
            I => \N__42327\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__42331\,
            I => \N__42324\
        );

    \I__9523\ : InMux
    port map (
            O => \N__42330\,
            I => \N__42321\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__42327\,
            I => \N__42318\
        );

    \I__9521\ : Span4Mux_v
    port map (
            O => \N__42324\,
            I => \N__42315\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__42321\,
            I => \N__42312\
        );

    \I__9519\ : Span4Mux_v
    port map (
            O => \N__42318\,
            I => \N__42308\
        );

    \I__9518\ : Span4Mux_v
    port map (
            O => \N__42315\,
            I => \N__42303\
        );

    \I__9517\ : Span4Mux_h
    port map (
            O => \N__42312\,
            I => \N__42303\
        );

    \I__9516\ : InMux
    port map (
            O => \N__42311\,
            I => \N__42300\
        );

    \I__9515\ : Odrv4
    port map (
            O => \N__42308\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__9514\ : Odrv4
    port map (
            O => \N__42303\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__42300\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__9512\ : InMux
    port map (
            O => \N__42293\,
            I => \N__42288\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42292\,
            I => \N__42285\
        );

    \I__9510\ : InMux
    port map (
            O => \N__42291\,
            I => \N__42282\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__42288\,
            I => \N__42279\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__42285\,
            I => \N__42276\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__42282\,
            I => \N__42271\
        );

    \I__9506\ : Span4Mux_v
    port map (
            O => \N__42279\,
            I => \N__42271\
        );

    \I__9505\ : Odrv4
    port map (
            O => \N__42276\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9504\ : Odrv4
    port map (
            O => \N__42271\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9503\ : CascadeMux
    port map (
            O => \N__42266\,
            I => \N__42263\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42263\,
            I => \N__42260\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__42260\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__9500\ : InMux
    port map (
            O => \N__42257\,
            I => \N__42242\
        );

    \I__9499\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42235\
        );

    \I__9498\ : InMux
    port map (
            O => \N__42255\,
            I => \N__42232\
        );

    \I__9497\ : InMux
    port map (
            O => \N__42254\,
            I => \N__42221\
        );

    \I__9496\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42221\
        );

    \I__9495\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42221\
        );

    \I__9494\ : InMux
    port map (
            O => \N__42251\,
            I => \N__42221\
        );

    \I__9493\ : InMux
    port map (
            O => \N__42250\,
            I => \N__42221\
        );

    \I__9492\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42205\
        );

    \I__9491\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42205\
        );

    \I__9490\ : InMux
    port map (
            O => \N__42247\,
            I => \N__42205\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42246\,
            I => \N__42205\
        );

    \I__9488\ : InMux
    port map (
            O => \N__42245\,
            I => \N__42205\
        );

    \I__9487\ : LocalMux
    port map (
            O => \N__42242\,
            I => \N__42202\
        );

    \I__9486\ : InMux
    port map (
            O => \N__42241\,
            I => \N__42193\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42240\,
            I => \N__42193\
        );

    \I__9484\ : InMux
    port map (
            O => \N__42239\,
            I => \N__42193\
        );

    \I__9483\ : InMux
    port map (
            O => \N__42238\,
            I => \N__42193\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__42235\,
            I => \N__42185\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__42232\,
            I => \N__42185\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__42221\,
            I => \N__42182\
        );

    \I__9479\ : InMux
    port map (
            O => \N__42220\,
            I => \N__42179\
        );

    \I__9478\ : InMux
    port map (
            O => \N__42219\,
            I => \N__42174\
        );

    \I__9477\ : InMux
    port map (
            O => \N__42218\,
            I => \N__42174\
        );

    \I__9476\ : InMux
    port map (
            O => \N__42217\,
            I => \N__42169\
        );

    \I__9475\ : InMux
    port map (
            O => \N__42216\,
            I => \N__42169\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__42205\,
            I => \N__42162\
        );

    \I__9473\ : Span4Mux_v
    port map (
            O => \N__42202\,
            I => \N__42162\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__42193\,
            I => \N__42162\
        );

    \I__9471\ : InMux
    port map (
            O => \N__42192\,
            I => \N__42159\
        );

    \I__9470\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42156\
        );

    \I__9469\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42153\
        );

    \I__9468\ : Span4Mux_v
    port map (
            O => \N__42185\,
            I => \N__42148\
        );

    \I__9467\ : Span4Mux_h
    port map (
            O => \N__42182\,
            I => \N__42148\
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__42179\,
            I => \N__42141\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__42174\,
            I => \N__42141\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__42169\,
            I => \N__42141\
        );

    \I__9463\ : Span4Mux_h
    port map (
            O => \N__42162\,
            I => \N__42138\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__42159\,
            I => \N__42133\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__42156\,
            I => \N__42133\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__42153\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9459\ : Odrv4
    port map (
            O => \N__42148\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9458\ : Odrv4
    port map (
            O => \N__42141\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9457\ : Odrv4
    port map (
            O => \N__42138\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9456\ : Odrv12
    port map (
            O => \N__42133\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__9455\ : CascadeMux
    port map (
            O => \N__42122\,
            I => \N__42118\
        );

    \I__9454\ : InMux
    port map (
            O => \N__42121\,
            I => \N__42115\
        );

    \I__9453\ : InMux
    port map (
            O => \N__42118\,
            I => \N__42112\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__42115\,
            I => \N__42108\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__42112\,
            I => \N__42105\
        );

    \I__9450\ : InMux
    port map (
            O => \N__42111\,
            I => \N__42102\
        );

    \I__9449\ : Span4Mux_v
    port map (
            O => \N__42108\,
            I => \N__42096\
        );

    \I__9448\ : Span4Mux_h
    port map (
            O => \N__42105\,
            I => \N__42096\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__42102\,
            I => \N__42093\
        );

    \I__9446\ : InMux
    port map (
            O => \N__42101\,
            I => \N__42090\
        );

    \I__9445\ : Odrv4
    port map (
            O => \N__42096\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9444\ : Odrv12
    port map (
            O => \N__42093\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__42090\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9442\ : InMux
    port map (
            O => \N__42083\,
            I => \N__42078\
        );

    \I__9441\ : InMux
    port map (
            O => \N__42082\,
            I => \N__42075\
        );

    \I__9440\ : CascadeMux
    port map (
            O => \N__42081\,
            I => \N__42072\
        );

    \I__9439\ : LocalMux
    port map (
            O => \N__42078\,
            I => \N__42067\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__42075\,
            I => \N__42067\
        );

    \I__9437\ : InMux
    port map (
            O => \N__42072\,
            I => \N__42064\
        );

    \I__9436\ : Span4Mux_v
    port map (
            O => \N__42067\,
            I => \N__42061\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__42064\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9434\ : Odrv4
    port map (
            O => \N__42061\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9433\ : CascadeMux
    port map (
            O => \N__42056\,
            I => \N__42053\
        );

    \I__9432\ : InMux
    port map (
            O => \N__42053\,
            I => \N__42050\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__42050\,
            I => \N__42047\
        );

    \I__9430\ : Odrv4
    port map (
            O => \N__42047\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__9429\ : InMux
    port map (
            O => \N__42044\,
            I => \N__42040\
        );

    \I__9428\ : InMux
    port map (
            O => \N__42043\,
            I => \N__42035\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__42040\,
            I => \N__42032\
        );

    \I__9426\ : InMux
    port map (
            O => \N__42039\,
            I => \N__42027\
        );

    \I__9425\ : InMux
    port map (
            O => \N__42038\,
            I => \N__42027\
        );

    \I__9424\ : LocalMux
    port map (
            O => \N__42035\,
            I => \N__42024\
        );

    \I__9423\ : Span4Mux_v
    port map (
            O => \N__42032\,
            I => \N__42019\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__42027\,
            I => \N__42019\
        );

    \I__9421\ : Odrv4
    port map (
            O => \N__42024\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9420\ : Odrv4
    port map (
            O => \N__42019\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9419\ : InMux
    port map (
            O => \N__42014\,
            I => \N__42011\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__42011\,
            I => \N__42007\
        );

    \I__9417\ : InMux
    port map (
            O => \N__42010\,
            I => \N__42004\
        );

    \I__9416\ : Span4Mux_h
    port map (
            O => \N__42007\,
            I => \N__42000\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__42004\,
            I => \N__41997\
        );

    \I__9414\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41994\
        );

    \I__9413\ : Odrv4
    port map (
            O => \N__42000\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__9412\ : Odrv4
    port map (
            O => \N__41997\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__41994\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__9410\ : CascadeMux
    port map (
            O => \N__41987\,
            I => \N__41983\
        );

    \I__9409\ : InMux
    port map (
            O => \N__41986\,
            I => \N__41979\
        );

    \I__9408\ : InMux
    port map (
            O => \N__41983\,
            I => \N__41976\
        );

    \I__9407\ : InMux
    port map (
            O => \N__41982\,
            I => \N__41973\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__41979\,
            I => \N__41969\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__41976\,
            I => \N__41966\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__41973\,
            I => \N__41963\
        );

    \I__9403\ : InMux
    port map (
            O => \N__41972\,
            I => \N__41959\
        );

    \I__9402\ : Span4Mux_v
    port map (
            O => \N__41969\,
            I => \N__41956\
        );

    \I__9401\ : Span4Mux_h
    port map (
            O => \N__41966\,
            I => \N__41953\
        );

    \I__9400\ : Span4Mux_h
    port map (
            O => \N__41963\,
            I => \N__41950\
        );

    \I__9399\ : InMux
    port map (
            O => \N__41962\,
            I => \N__41947\
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__41959\,
            I => \N__41943\
        );

    \I__9397\ : Span4Mux_h
    port map (
            O => \N__41956\,
            I => \N__41938\
        );

    \I__9396\ : Span4Mux_v
    port map (
            O => \N__41953\,
            I => \N__41938\
        );

    \I__9395\ : Span4Mux_v
    port map (
            O => \N__41950\,
            I => \N__41935\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__41947\,
            I => \N__41932\
        );

    \I__9393\ : InMux
    port map (
            O => \N__41946\,
            I => \N__41929\
        );

    \I__9392\ : Span4Mux_v
    port map (
            O => \N__41943\,
            I => \N__41926\
        );

    \I__9391\ : Span4Mux_v
    port map (
            O => \N__41938\,
            I => \N__41923\
        );

    \I__9390\ : Sp12to4
    port map (
            O => \N__41935\,
            I => \N__41918\
        );

    \I__9389\ : Span12Mux_h
    port map (
            O => \N__41932\,
            I => \N__41918\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__41929\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__9387\ : Odrv4
    port map (
            O => \N__41926\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__9386\ : Odrv4
    port map (
            O => \N__41923\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__9385\ : Odrv12
    port map (
            O => \N__41918\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__9384\ : IoInMux
    port map (
            O => \N__41909\,
            I => \N__41906\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__41906\,
            I => \N__41903\
        );

    \I__9382\ : IoSpan4Mux
    port map (
            O => \N__41903\,
            I => \N__41900\
        );

    \I__9381\ : Sp12to4
    port map (
            O => \N__41900\,
            I => \N__41896\
        );

    \I__9380\ : InMux
    port map (
            O => \N__41899\,
            I => \N__41893\
        );

    \I__9379\ : Odrv12
    port map (
            O => \N__41896\,
            I => \T01_c\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__41893\,
            I => \T01_c\
        );

    \I__9377\ : InMux
    port map (
            O => \N__41888\,
            I => \N__41884\
        );

    \I__9376\ : InMux
    port map (
            O => \N__41887\,
            I => \N__41881\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__41884\,
            I => \N__41876\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__41881\,
            I => \N__41873\
        );

    \I__9373\ : InMux
    port map (
            O => \N__41880\,
            I => \N__41868\
        );

    \I__9372\ : InMux
    port map (
            O => \N__41879\,
            I => \N__41868\
        );

    \I__9371\ : Span4Mux_h
    port map (
            O => \N__41876\,
            I => \N__41865\
        );

    \I__9370\ : Odrv12
    port map (
            O => \N__41873\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__41868\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__9368\ : Odrv4
    port map (
            O => \N__41865\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__9367\ : InMux
    port map (
            O => \N__41858\,
            I => \N__41854\
        );

    \I__9366\ : InMux
    port map (
            O => \N__41857\,
            I => \N__41851\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__41854\,
            I => \N__41847\
        );

    \I__9364\ : LocalMux
    port map (
            O => \N__41851\,
            I => \N__41843\
        );

    \I__9363\ : InMux
    port map (
            O => \N__41850\,
            I => \N__41840\
        );

    \I__9362\ : Span4Mux_v
    port map (
            O => \N__41847\,
            I => \N__41837\
        );

    \I__9361\ : InMux
    port map (
            O => \N__41846\,
            I => \N__41834\
        );

    \I__9360\ : Span4Mux_h
    port map (
            O => \N__41843\,
            I => \N__41831\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__41840\,
            I => \N__41827\
        );

    \I__9358\ : Sp12to4
    port map (
            O => \N__41837\,
            I => \N__41822\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__41834\,
            I => \N__41822\
        );

    \I__9356\ : Span4Mux_h
    port map (
            O => \N__41831\,
            I => \N__41819\
        );

    \I__9355\ : InMux
    port map (
            O => \N__41830\,
            I => \N__41816\
        );

    \I__9354\ : Span4Mux_v
    port map (
            O => \N__41827\,
            I => \N__41813\
        );

    \I__9353\ : Odrv12
    port map (
            O => \N__41822\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__9352\ : Odrv4
    port map (
            O => \N__41819\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__41816\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__9350\ : Odrv4
    port map (
            O => \N__41813\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__9349\ : IoInMux
    port map (
            O => \N__41804\,
            I => \N__41801\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__41801\,
            I => \N__41798\
        );

    \I__9347\ : Span4Mux_s3_v
    port map (
            O => \N__41798\,
            I => \N__41794\
        );

    \I__9346\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41791\
        );

    \I__9345\ : Odrv4
    port map (
            O => \N__41794\,
            I => \T12_c\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__41791\,
            I => \T12_c\
        );

    \I__9343\ : InMux
    port map (
            O => \N__41786\,
            I => \N__41782\
        );

    \I__9342\ : InMux
    port map (
            O => \N__41785\,
            I => \N__41779\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__41782\,
            I => \N__41775\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__41779\,
            I => \N__41772\
        );

    \I__9339\ : InMux
    port map (
            O => \N__41778\,
            I => \N__41769\
        );

    \I__9338\ : Span4Mux_v
    port map (
            O => \N__41775\,
            I => \N__41765\
        );

    \I__9337\ : Span4Mux_v
    port map (
            O => \N__41772\,
            I => \N__41760\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__41769\,
            I => \N__41760\
        );

    \I__9335\ : InMux
    port map (
            O => \N__41768\,
            I => \N__41757\
        );

    \I__9334\ : Odrv4
    port map (
            O => \N__41765\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9333\ : Odrv4
    port map (
            O => \N__41760\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__41757\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9331\ : CascadeMux
    port map (
            O => \N__41750\,
            I => \N__41746\
        );

    \I__9330\ : CascadeMux
    port map (
            O => \N__41749\,
            I => \N__41743\
        );

    \I__9329\ : InMux
    port map (
            O => \N__41746\,
            I => \N__41740\
        );

    \I__9328\ : InMux
    port map (
            O => \N__41743\,
            I => \N__41737\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__41740\,
            I => \N__41734\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__41737\,
            I => \N__41730\
        );

    \I__9325\ : Span4Mux_h
    port map (
            O => \N__41734\,
            I => \N__41727\
        );

    \I__9324\ : InMux
    port map (
            O => \N__41733\,
            I => \N__41724\
        );

    \I__9323\ : Odrv4
    port map (
            O => \N__41730\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9322\ : Odrv4
    port map (
            O => \N__41727\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__41724\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9320\ : InMux
    port map (
            O => \N__41717\,
            I => \N__41712\
        );

    \I__9319\ : InMux
    port map (
            O => \N__41716\,
            I => \N__41705\
        );

    \I__9318\ : InMux
    port map (
            O => \N__41715\,
            I => \N__41705\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__41712\,
            I => \N__41685\
        );

    \I__9316\ : InMux
    port map (
            O => \N__41711\,
            I => \N__41682\
        );

    \I__9315\ : InMux
    port map (
            O => \N__41710\,
            I => \N__41679\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__41705\,
            I => \N__41676\
        );

    \I__9313\ : InMux
    port map (
            O => \N__41704\,
            I => \N__41671\
        );

    \I__9312\ : InMux
    port map (
            O => \N__41703\,
            I => \N__41671\
        );

    \I__9311\ : InMux
    port map (
            O => \N__41702\,
            I => \N__41668\
        );

    \I__9310\ : InMux
    port map (
            O => \N__41701\,
            I => \N__41663\
        );

    \I__9309\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41663\
        );

    \I__9308\ : InMux
    port map (
            O => \N__41699\,
            I => \N__41656\
        );

    \I__9307\ : InMux
    port map (
            O => \N__41698\,
            I => \N__41656\
        );

    \I__9306\ : InMux
    port map (
            O => \N__41697\,
            I => \N__41656\
        );

    \I__9305\ : InMux
    port map (
            O => \N__41696\,
            I => \N__41649\
        );

    \I__9304\ : InMux
    port map (
            O => \N__41695\,
            I => \N__41649\
        );

    \I__9303\ : InMux
    port map (
            O => \N__41694\,
            I => \N__41649\
        );

    \I__9302\ : InMux
    port map (
            O => \N__41693\,
            I => \N__41638\
        );

    \I__9301\ : InMux
    port map (
            O => \N__41692\,
            I => \N__41638\
        );

    \I__9300\ : InMux
    port map (
            O => \N__41691\,
            I => \N__41638\
        );

    \I__9299\ : InMux
    port map (
            O => \N__41690\,
            I => \N__41638\
        );

    \I__9298\ : InMux
    port map (
            O => \N__41689\,
            I => \N__41638\
        );

    \I__9297\ : InMux
    port map (
            O => \N__41688\,
            I => \N__41635\
        );

    \I__9296\ : Span12Mux_v
    port map (
            O => \N__41685\,
            I => \N__41630\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__41682\,
            I => \N__41630\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__41679\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__9293\ : Odrv4
    port map (
            O => \N__41676\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__41671\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__41668\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__41663\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__41656\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__41649\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__41638\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__41635\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__9285\ : Odrv12
    port map (
            O => \N__41630\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__9284\ : InMux
    port map (
            O => \N__41609\,
            I => \N__41606\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__41606\,
            I => \N__41602\
        );

    \I__9282\ : CascadeMux
    port map (
            O => \N__41605\,
            I => \N__41598\
        );

    \I__9281\ : Span12Mux_v
    port map (
            O => \N__41602\,
            I => \N__41595\
        );

    \I__9280\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41590\
        );

    \I__9279\ : InMux
    port map (
            O => \N__41598\,
            I => \N__41590\
        );

    \I__9278\ : Span12Mux_h
    port map (
            O => \N__41595\,
            I => \N__41587\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__41590\,
            I => \N__41584\
        );

    \I__9276\ : Odrv12
    port map (
            O => \N__41587\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__9275\ : Odrv12
    port map (
            O => \N__41584\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__41579\,
            I => \N__41576\
        );

    \I__9273\ : InMux
    port map (
            O => \N__41576\,
            I => \N__41570\
        );

    \I__9272\ : InMux
    port map (
            O => \N__41575\,
            I => \N__41558\
        );

    \I__9271\ : InMux
    port map (
            O => \N__41574\,
            I => \N__41558\
        );

    \I__9270\ : CascadeMux
    port map (
            O => \N__41573\,
            I => \N__41555\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__41570\,
            I => \N__41552\
        );

    \I__9268\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41546\
        );

    \I__9267\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41541\
        );

    \I__9266\ : InMux
    port map (
            O => \N__41567\,
            I => \N__41534\
        );

    \I__9265\ : InMux
    port map (
            O => \N__41566\,
            I => \N__41534\
        );

    \I__9264\ : InMux
    port map (
            O => \N__41565\,
            I => \N__41534\
        );

    \I__9263\ : CascadeMux
    port map (
            O => \N__41564\,
            I => \N__41531\
        );

    \I__9262\ : CascadeMux
    port map (
            O => \N__41563\,
            I => \N__41527\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__41558\,
            I => \N__41524\
        );

    \I__9260\ : InMux
    port map (
            O => \N__41555\,
            I => \N__41515\
        );

    \I__9259\ : Span4Mux_h
    port map (
            O => \N__41552\,
            I => \N__41512\
        );

    \I__9258\ : CascadeMux
    port map (
            O => \N__41551\,
            I => \N__41508\
        );

    \I__9257\ : CascadeMux
    port map (
            O => \N__41550\,
            I => \N__41505\
        );

    \I__9256\ : CascadeMux
    port map (
            O => \N__41549\,
            I => \N__41501\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__41546\,
            I => \N__41493\
        );

    \I__9254\ : InMux
    port map (
            O => \N__41545\,
            I => \N__41490\
        );

    \I__9253\ : InMux
    port map (
            O => \N__41544\,
            I => \N__41487\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__41541\,
            I => \N__41484\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__41534\,
            I => \N__41481\
        );

    \I__9250\ : InMux
    port map (
            O => \N__41531\,
            I => \N__41478\
        );

    \I__9249\ : InMux
    port map (
            O => \N__41530\,
            I => \N__41475\
        );

    \I__9248\ : InMux
    port map (
            O => \N__41527\,
            I => \N__41472\
        );

    \I__9247\ : Span4Mux_h
    port map (
            O => \N__41524\,
            I => \N__41469\
        );

    \I__9246\ : InMux
    port map (
            O => \N__41523\,
            I => \N__41464\
        );

    \I__9245\ : InMux
    port map (
            O => \N__41522\,
            I => \N__41464\
        );

    \I__9244\ : InMux
    port map (
            O => \N__41521\,
            I => \N__41461\
        );

    \I__9243\ : InMux
    port map (
            O => \N__41520\,
            I => \N__41454\
        );

    \I__9242\ : InMux
    port map (
            O => \N__41519\,
            I => \N__41454\
        );

    \I__9241\ : InMux
    port map (
            O => \N__41518\,
            I => \N__41454\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__41515\,
            I => \N__41449\
        );

    \I__9239\ : Span4Mux_h
    port map (
            O => \N__41512\,
            I => \N__41449\
        );

    \I__9238\ : InMux
    port map (
            O => \N__41511\,
            I => \N__41444\
        );

    \I__9237\ : InMux
    port map (
            O => \N__41508\,
            I => \N__41444\
        );

    \I__9236\ : InMux
    port map (
            O => \N__41505\,
            I => \N__41441\
        );

    \I__9235\ : InMux
    port map (
            O => \N__41504\,
            I => \N__41434\
        );

    \I__9234\ : InMux
    port map (
            O => \N__41501\,
            I => \N__41434\
        );

    \I__9233\ : InMux
    port map (
            O => \N__41500\,
            I => \N__41434\
        );

    \I__9232\ : InMux
    port map (
            O => \N__41499\,
            I => \N__41425\
        );

    \I__9231\ : InMux
    port map (
            O => \N__41498\,
            I => \N__41425\
        );

    \I__9230\ : InMux
    port map (
            O => \N__41497\,
            I => \N__41425\
        );

    \I__9229\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41425\
        );

    \I__9228\ : Span4Mux_v
    port map (
            O => \N__41493\,
            I => \N__41416\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__41490\,
            I => \N__41416\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__41487\,
            I => \N__41416\
        );

    \I__9225\ : Span4Mux_v
    port map (
            O => \N__41484\,
            I => \N__41416\
        );

    \I__9224\ : Odrv12
    port map (
            O => \N__41481\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__41478\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__41475\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__41472\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9220\ : Odrv4
    port map (
            O => \N__41469\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__41464\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__41461\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__41454\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9216\ : Odrv4
    port map (
            O => \N__41449\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__41444\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__41441\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__41434\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__41425\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9211\ : Odrv4
    port map (
            O => \N__41416\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__9210\ : InMux
    port map (
            O => \N__41387\,
            I => \N__41383\
        );

    \I__9209\ : InMux
    port map (
            O => \N__41386\,
            I => \N__41380\
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__41383\,
            I => \N__41377\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__41380\,
            I => \N__41374\
        );

    \I__9206\ : Span4Mux_v
    port map (
            O => \N__41377\,
            I => \N__41370\
        );

    \I__9205\ : Span4Mux_v
    port map (
            O => \N__41374\,
            I => \N__41367\
        );

    \I__9204\ : InMux
    port map (
            O => \N__41373\,
            I => \N__41364\
        );

    \I__9203\ : Sp12to4
    port map (
            O => \N__41370\,
            I => \N__41359\
        );

    \I__9202\ : Sp12to4
    port map (
            O => \N__41367\,
            I => \N__41359\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__41364\,
            I => \elapsed_time_ns_1_RNI81DJ11_0_2\
        );

    \I__9200\ : Odrv12
    port map (
            O => \N__41359\,
            I => \elapsed_time_ns_1_RNI81DJ11_0_2\
        );

    \I__9199\ : CascadeMux
    port map (
            O => \N__41354\,
            I => \N__41350\
        );

    \I__9198\ : CascadeMux
    port map (
            O => \N__41353\,
            I => \N__41347\
        );

    \I__9197\ : InMux
    port map (
            O => \N__41350\,
            I => \N__41344\
        );

    \I__9196\ : InMux
    port map (
            O => \N__41347\,
            I => \N__41341\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__41344\,
            I => \N__41337\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__41341\,
            I => \N__41334\
        );

    \I__9193\ : InMux
    port map (
            O => \N__41340\,
            I => \N__41331\
        );

    \I__9192\ : Span4Mux_v
    port map (
            O => \N__41337\,
            I => \N__41328\
        );

    \I__9191\ : Span4Mux_v
    port map (
            O => \N__41334\,
            I => \N__41325\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__41331\,
            I => \N__41322\
        );

    \I__9189\ : Span4Mux_v
    port map (
            O => \N__41328\,
            I => \N__41318\
        );

    \I__9188\ : Span4Mux_v
    port map (
            O => \N__41325\,
            I => \N__41313\
        );

    \I__9187\ : Span4Mux_h
    port map (
            O => \N__41322\,
            I => \N__41313\
        );

    \I__9186\ : InMux
    port map (
            O => \N__41321\,
            I => \N__41310\
        );

    \I__9185\ : Odrv4
    port map (
            O => \N__41318\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__9184\ : Odrv4
    port map (
            O => \N__41313\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__41310\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__9182\ : InMux
    port map (
            O => \N__41303\,
            I => \N__41299\
        );

    \I__9181\ : InMux
    port map (
            O => \N__41302\,
            I => \N__41296\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__41299\,
            I => \N__41293\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__41296\,
            I => \N__41289\
        );

    \I__9178\ : Span4Mux_h
    port map (
            O => \N__41293\,
            I => \N__41286\
        );

    \I__9177\ : InMux
    port map (
            O => \N__41292\,
            I => \N__41283\
        );

    \I__9176\ : Odrv12
    port map (
            O => \N__41289\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9175\ : Odrv4
    port map (
            O => \N__41286\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__41283\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9173\ : InMux
    port map (
            O => \N__41276\,
            I => \N__41273\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__41273\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__9171\ : CascadeMux
    port map (
            O => \N__41270\,
            I => \N__41267\
        );

    \I__9170\ : InMux
    port map (
            O => \N__41267\,
            I => \N__41264\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__41264\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__9168\ : InMux
    port map (
            O => \N__41261\,
            I => \N__41257\
        );

    \I__9167\ : CascadeMux
    port map (
            O => \N__41260\,
            I => \N__41254\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__41257\,
            I => \N__41250\
        );

    \I__9165\ : InMux
    port map (
            O => \N__41254\,
            I => \N__41247\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41253\,
            I => \N__41244\
        );

    \I__9163\ : Span4Mux_h
    port map (
            O => \N__41250\,
            I => \N__41241\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__41247\,
            I => \N__41236\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__41244\,
            I => \N__41236\
        );

    \I__9160\ : Odrv4
    port map (
            O => \N__41241\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9159\ : Odrv4
    port map (
            O => \N__41236\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9158\ : CascadeMux
    port map (
            O => \N__41231\,
            I => \N__41228\
        );

    \I__9157\ : InMux
    port map (
            O => \N__41228\,
            I => \N__41223\
        );

    \I__9156\ : InMux
    port map (
            O => \N__41227\,
            I => \N__41218\
        );

    \I__9155\ : InMux
    port map (
            O => \N__41226\,
            I => \N__41218\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__41223\,
            I => \N__41215\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__41218\,
            I => \N__41212\
        );

    \I__9152\ : Span4Mux_v
    port map (
            O => \N__41215\,
            I => \N__41206\
        );

    \I__9151\ : Span4Mux_h
    port map (
            O => \N__41212\,
            I => \N__41206\
        );

    \I__9150\ : InMux
    port map (
            O => \N__41211\,
            I => \N__41203\
        );

    \I__9149\ : Odrv4
    port map (
            O => \N__41206\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__41203\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__9147\ : InMux
    port map (
            O => \N__41198\,
            I => \N__41189\
        );

    \I__9146\ : InMux
    port map (
            O => \N__41197\,
            I => \N__41189\
        );

    \I__9145\ : InMux
    port map (
            O => \N__41196\,
            I => \N__41189\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__41189\,
            I => \N__41186\
        );

    \I__9143\ : Span4Mux_v
    port map (
            O => \N__41186\,
            I => \N__41183\
        );

    \I__9142\ : Span4Mux_v
    port map (
            O => \N__41183\,
            I => \N__41179\
        );

    \I__9141\ : InMux
    port map (
            O => \N__41182\,
            I => \N__41176\
        );

    \I__9140\ : Odrv4
    port map (
            O => \N__41179\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__41176\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__9138\ : CascadeMux
    port map (
            O => \N__41171\,
            I => \N__41168\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41168\,
            I => \N__41159\
        );

    \I__9136\ : InMux
    port map (
            O => \N__41167\,
            I => \N__41159\
        );

    \I__9135\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41159\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__41159\,
            I => \N__41156\
        );

    \I__9133\ : Span4Mux_h
    port map (
            O => \N__41156\,
            I => \N__41153\
        );

    \I__9132\ : Odrv4
    port map (
            O => \N__41153\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9131\ : CascadeMux
    port map (
            O => \N__41150\,
            I => \N__41147\
        );

    \I__9130\ : InMux
    port map (
            O => \N__41147\,
            I => \N__41144\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__41144\,
            I => \N__41141\
        );

    \I__9128\ : Odrv4
    port map (
            O => \N__41141\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__9127\ : InMux
    port map (
            O => \N__41138\,
            I => \N__41135\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__41135\,
            I => \N__41132\
        );

    \I__9125\ : Odrv4
    port map (
            O => \N__41132\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__9124\ : InMux
    port map (
            O => \N__41129\,
            I => \N__41126\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__41126\,
            I => \N__41123\
        );

    \I__9122\ : Span4Mux_h
    port map (
            O => \N__41123\,
            I => \N__41120\
        );

    \I__9121\ : Odrv4
    port map (
            O => \N__41120\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__9120\ : InMux
    port map (
            O => \N__41117\,
            I => \N__41108\
        );

    \I__9119\ : InMux
    port map (
            O => \N__41116\,
            I => \N__41108\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41115\,
            I => \N__41108\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__41108\,
            I => \N__41105\
        );

    \I__9116\ : Span4Mux_h
    port map (
            O => \N__41105\,
            I => \N__41102\
        );

    \I__9115\ : Span4Mux_v
    port map (
            O => \N__41102\,
            I => \N__41098\
        );

    \I__9114\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41095\
        );

    \I__9113\ : Odrv4
    port map (
            O => \N__41098\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__41095\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9111\ : CascadeMux
    port map (
            O => \N__41090\,
            I => \N__41087\
        );

    \I__9110\ : InMux
    port map (
            O => \N__41087\,
            I => \N__41078\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41086\,
            I => \N__41078\
        );

    \I__9108\ : InMux
    port map (
            O => \N__41085\,
            I => \N__41078\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__41078\,
            I => \N__41075\
        );

    \I__9106\ : Span4Mux_h
    port map (
            O => \N__41075\,
            I => \N__41072\
        );

    \I__9105\ : Odrv4
    port map (
            O => \N__41072\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9104\ : CascadeMux
    port map (
            O => \N__41069\,
            I => \N__41066\
        );

    \I__9103\ : InMux
    port map (
            O => \N__41066\,
            I => \N__41063\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__41063\,
            I => \N__41060\
        );

    \I__9101\ : Odrv4
    port map (
            O => \N__41060\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__9100\ : InMux
    port map (
            O => \N__41057\,
            I => \N__41054\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__41054\,
            I => \N__41049\
        );

    \I__9098\ : InMux
    port map (
            O => \N__41053\,
            I => \N__41046\
        );

    \I__9097\ : InMux
    port map (
            O => \N__41052\,
            I => \N__41043\
        );

    \I__9096\ : Span4Mux_h
    port map (
            O => \N__41049\,
            I => \N__41038\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__41046\,
            I => \N__41038\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41043\,
            I => \N__41035\
        );

    \I__9093\ : Span4Mux_v
    port map (
            O => \N__41038\,
            I => \N__41030\
        );

    \I__9092\ : Span4Mux_h
    port map (
            O => \N__41035\,
            I => \N__41030\
        );

    \I__9091\ : Span4Mux_v
    port map (
            O => \N__41030\,
            I => \N__41027\
        );

    \I__9090\ : Odrv4
    port map (
            O => \N__41027\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__9089\ : CEMux
    port map (
            O => \N__41024\,
            I => \N__40997\
        );

    \I__9088\ : CEMux
    port map (
            O => \N__41023\,
            I => \N__40997\
        );

    \I__9087\ : CEMux
    port map (
            O => \N__41022\,
            I => \N__40997\
        );

    \I__9086\ : CEMux
    port map (
            O => \N__41021\,
            I => \N__40997\
        );

    \I__9085\ : CEMux
    port map (
            O => \N__41020\,
            I => \N__40997\
        );

    \I__9084\ : CEMux
    port map (
            O => \N__41019\,
            I => \N__40997\
        );

    \I__9083\ : CEMux
    port map (
            O => \N__41018\,
            I => \N__40997\
        );

    \I__9082\ : CEMux
    port map (
            O => \N__41017\,
            I => \N__40997\
        );

    \I__9081\ : CEMux
    port map (
            O => \N__41016\,
            I => \N__40997\
        );

    \I__9080\ : GlobalMux
    port map (
            O => \N__40997\,
            I => \N__40994\
        );

    \I__9079\ : gio2CtrlBuf
    port map (
            O => \N__40994\,
            I => \current_shift_inst.timer_s1.N_166_i_g\
        );

    \I__9078\ : InMux
    port map (
            O => \N__40991\,
            I => \N__40988\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__40988\,
            I => \N__40985\
        );

    \I__9076\ : Span4Mux_h
    port map (
            O => \N__40985\,
            I => \N__40982\
        );

    \I__9075\ : Odrv4
    port map (
            O => \N__40982\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__9074\ : InMux
    port map (
            O => \N__40979\,
            I => \N__40976\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__40976\,
            I => \N__40973\
        );

    \I__9072\ : Odrv4
    port map (
            O => \N__40973\,
            I => \current_shift_inst.control_input_1_axb_6\
        );

    \I__9071\ : InMux
    port map (
            O => \N__40970\,
            I => \N__40967\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__40967\,
            I => \N__40964\
        );

    \I__9069\ : Span4Mux_v
    port map (
            O => \N__40964\,
            I => \N__40961\
        );

    \I__9068\ : Odrv4
    port map (
            O => \N__40961\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__9067\ : InMux
    port map (
            O => \N__40958\,
            I => \N__40955\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__40955\,
            I => \N__40952\
        );

    \I__9065\ : Odrv4
    port map (
            O => \N__40952\,
            I => \current_shift_inst.control_input_1_axb_8\
        );

    \I__9064\ : InMux
    port map (
            O => \N__40949\,
            I => \N__40946\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__40946\,
            I => \N__40943\
        );

    \I__9062\ : Span4Mux_v
    port map (
            O => \N__40943\,
            I => \N__40940\
        );

    \I__9061\ : Odrv4
    port map (
            O => \N__40940\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__9060\ : InMux
    port map (
            O => \N__40937\,
            I => \N__40922\
        );

    \I__9059\ : InMux
    port map (
            O => \N__40936\,
            I => \N__40913\
        );

    \I__9058\ : InMux
    port map (
            O => \N__40935\,
            I => \N__40913\
        );

    \I__9057\ : InMux
    port map (
            O => \N__40934\,
            I => \N__40913\
        );

    \I__9056\ : InMux
    port map (
            O => \N__40933\,
            I => \N__40913\
        );

    \I__9055\ : InMux
    port map (
            O => \N__40932\,
            I => \N__40902\
        );

    \I__9054\ : InMux
    port map (
            O => \N__40931\,
            I => \N__40902\
        );

    \I__9053\ : InMux
    port map (
            O => \N__40930\,
            I => \N__40902\
        );

    \I__9052\ : InMux
    port map (
            O => \N__40929\,
            I => \N__40902\
        );

    \I__9051\ : InMux
    port map (
            O => \N__40928\,
            I => \N__40902\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40927\,
            I => \N__40895\
        );

    \I__9049\ : InMux
    port map (
            O => \N__40926\,
            I => \N__40895\
        );

    \I__9048\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40895\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__40922\,
            I => \N__40888\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__40913\,
            I => \N__40888\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__40902\,
            I => \N__40888\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__40895\,
            I => \N__40885\
        );

    \I__9043\ : Span4Mux_v
    port map (
            O => \N__40888\,
            I => \N__40882\
        );

    \I__9042\ : Odrv4
    port map (
            O => \N__40885\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9041\ : Odrv4
    port map (
            O => \N__40882\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__9040\ : InMux
    port map (
            O => \N__40877\,
            I => \N__40874\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__40874\,
            I => \N__40871\
        );

    \I__9038\ : Odrv4
    port map (
            O => \N__40871\,
            I => \current_shift_inst.control_input_1_axb_9\
        );

    \I__9037\ : InMux
    port map (
            O => \N__40868\,
            I => \N__40864\
        );

    \I__9036\ : InMux
    port map (
            O => \N__40867\,
            I => \N__40861\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__40864\,
            I => \N__40858\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__40861\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__9033\ : Odrv4
    port map (
            O => \N__40858\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__9032\ : InMux
    port map (
            O => \N__40853\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__9031\ : InMux
    port map (
            O => \N__40850\,
            I => \N__40847\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__40847\,
            I => \N__40843\
        );

    \I__9029\ : InMux
    port map (
            O => \N__40846\,
            I => \N__40840\
        );

    \I__9028\ : Span4Mux_h
    port map (
            O => \N__40843\,
            I => \N__40837\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__40840\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__9026\ : Odrv4
    port map (
            O => \N__40837\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__9025\ : InMux
    port map (
            O => \N__40832\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__9024\ : InMux
    port map (
            O => \N__40829\,
            I => \N__40825\
        );

    \I__9023\ : InMux
    port map (
            O => \N__40828\,
            I => \N__40822\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__40825\,
            I => \N__40819\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__40822\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9020\ : Odrv12
    port map (
            O => \N__40819\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9019\ : InMux
    port map (
            O => \N__40814\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__9018\ : InMux
    port map (
            O => \N__40811\,
            I => \N__40807\
        );

    \I__9017\ : InMux
    port map (
            O => \N__40810\,
            I => \N__40804\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__40807\,
            I => \N__40801\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__40804\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9014\ : Odrv4
    port map (
            O => \N__40801\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9013\ : InMux
    port map (
            O => \N__40796\,
            I => \bfn_17_16_0_\
        );

    \I__9012\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40789\
        );

    \I__9011\ : InMux
    port map (
            O => \N__40792\,
            I => \N__40786\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__40789\,
            I => \N__40783\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__40786\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9008\ : Odrv4
    port map (
            O => \N__40783\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9007\ : InMux
    port map (
            O => \N__40778\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__9006\ : InMux
    port map (
            O => \N__40775\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__9005\ : InMux
    port map (
            O => \N__40772\,
            I => \N__40768\
        );

    \I__9004\ : InMux
    port map (
            O => \N__40771\,
            I => \N__40765\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__40768\,
            I => \N__40762\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__40765\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9001\ : Odrv4
    port map (
            O => \N__40762\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9000\ : CascadeMux
    port map (
            O => \N__40757\,
            I => \N__40754\
        );

    \I__8999\ : InMux
    port map (
            O => \N__40754\,
            I => \N__40751\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__40751\,
            I => \N__40748\
        );

    \I__8997\ : Odrv4
    port map (
            O => \N__40748\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__8996\ : InMux
    port map (
            O => \N__40745\,
            I => \N__40741\
        );

    \I__8995\ : InMux
    port map (
            O => \N__40744\,
            I => \N__40738\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__40741\,
            I => \N__40735\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__40738\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8992\ : Odrv4
    port map (
            O => \N__40735\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8991\ : InMux
    port map (
            O => \N__40730\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__8990\ : InMux
    port map (
            O => \N__40727\,
            I => \N__40723\
        );

    \I__8989\ : InMux
    port map (
            O => \N__40726\,
            I => \N__40720\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__40723\,
            I => \N__40717\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__40720\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8986\ : Odrv4
    port map (
            O => \N__40717\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8985\ : InMux
    port map (
            O => \N__40712\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__8984\ : InMux
    port map (
            O => \N__40709\,
            I => \N__40705\
        );

    \I__8983\ : InMux
    port map (
            O => \N__40708\,
            I => \N__40702\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__40705\,
            I => \N__40699\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__40702\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8980\ : Odrv12
    port map (
            O => \N__40699\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8979\ : InMux
    port map (
            O => \N__40694\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__8978\ : InMux
    port map (
            O => \N__40691\,
            I => \N__40687\
        );

    \I__8977\ : InMux
    port map (
            O => \N__40690\,
            I => \N__40684\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__40687\,
            I => \N__40681\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__40684\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8974\ : Odrv12
    port map (
            O => \N__40681\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8973\ : InMux
    port map (
            O => \N__40676\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__8972\ : InMux
    port map (
            O => \N__40673\,
            I => \N__40669\
        );

    \I__8971\ : InMux
    port map (
            O => \N__40672\,
            I => \N__40666\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__40669\,
            I => \N__40663\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__40666\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8968\ : Odrv4
    port map (
            O => \N__40663\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8967\ : InMux
    port map (
            O => \N__40658\,
            I => \bfn_17_15_0_\
        );

    \I__8966\ : InMux
    port map (
            O => \N__40655\,
            I => \N__40651\
        );

    \I__8965\ : InMux
    port map (
            O => \N__40654\,
            I => \N__40648\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__40651\,
            I => \N__40645\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__40648\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8962\ : Odrv4
    port map (
            O => \N__40645\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8961\ : InMux
    port map (
            O => \N__40640\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__8960\ : InMux
    port map (
            O => \N__40637\,
            I => \N__40633\
        );

    \I__8959\ : InMux
    port map (
            O => \N__40636\,
            I => \N__40630\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__40633\,
            I => \N__40627\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__40630\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8956\ : Odrv4
    port map (
            O => \N__40627\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8955\ : InMux
    port map (
            O => \N__40622\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__8954\ : InMux
    port map (
            O => \N__40619\,
            I => \N__40615\
        );

    \I__8953\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40612\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__40615\,
            I => \N__40609\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__40612\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8950\ : Odrv4
    port map (
            O => \N__40609\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8949\ : InMux
    port map (
            O => \N__40604\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__8948\ : InMux
    port map (
            O => \N__40601\,
            I => \N__40597\
        );

    \I__8947\ : InMux
    port map (
            O => \N__40600\,
            I => \N__40594\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__40597\,
            I => \N__40591\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__40594\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8944\ : Odrv4
    port map (
            O => \N__40591\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8943\ : InMux
    port map (
            O => \N__40586\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__8942\ : InMux
    port map (
            O => \N__40583\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_19\
        );

    \I__8941\ : InMux
    port map (
            O => \N__40580\,
            I => \N__40577\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__40577\,
            I => \N__40573\
        );

    \I__8939\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40570\
        );

    \I__8938\ : Span4Mux_s1_v
    port map (
            O => \N__40573\,
            I => \N__40565\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__40570\,
            I => \N__40565\
        );

    \I__8936\ : Span4Mux_v
    port map (
            O => \N__40565\,
            I => \N__40561\
        );

    \I__8935\ : InMux
    port map (
            O => \N__40564\,
            I => \N__40558\
        );

    \I__8934\ : Span4Mux_h
    port map (
            O => \N__40561\,
            I => \N__40555\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__40558\,
            I => \N__40552\
        );

    \I__8932\ : Sp12to4
    port map (
            O => \N__40555\,
            I => \N__40548\
        );

    \I__8931\ : Span4Mux_v
    port map (
            O => \N__40552\,
            I => \N__40545\
        );

    \I__8930\ : InMux
    port map (
            O => \N__40551\,
            I => \N__40542\
        );

    \I__8929\ : Span12Mux_v
    port map (
            O => \N__40548\,
            I => \N__40539\
        );

    \I__8928\ : Span4Mux_h
    port map (
            O => \N__40545\,
            I => \N__40534\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__40542\,
            I => \N__40534\
        );

    \I__8926\ : Span12Mux_v
    port map (
            O => \N__40539\,
            I => \N__40531\
        );

    \I__8925\ : Span4Mux_v
    port map (
            O => \N__40534\,
            I => \N__40528\
        );

    \I__8924\ : Span12Mux_h
    port map (
            O => \N__40531\,
            I => \N__40525\
        );

    \I__8923\ : Sp12to4
    port map (
            O => \N__40528\,
            I => \N__40522\
        );

    \I__8922\ : Odrv12
    port map (
            O => \N__40525\,
            I => start_stop_c
        );

    \I__8921\ : Odrv12
    port map (
            O => \N__40522\,
            I => start_stop_c
        );

    \I__8920\ : InMux
    port map (
            O => \N__40517\,
            I => \N__40514\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__40514\,
            I => \N__40510\
        );

    \I__8918\ : InMux
    port map (
            O => \N__40513\,
            I => \N__40507\
        );

    \I__8917\ : Span4Mux_v
    port map (
            O => \N__40510\,
            I => \N__40502\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__40507\,
            I => \N__40502\
        );

    \I__8915\ : Span4Mux_h
    port map (
            O => \N__40502\,
            I => \N__40499\
        );

    \I__8914\ : Odrv4
    port map (
            O => \N__40499\,
            I => state_ns_i_a3_1
        );

    \I__8913\ : InMux
    port map (
            O => \N__40496\,
            I => \N__40493\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__40493\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__8911\ : InMux
    port map (
            O => \N__40490\,
            I => \N__40486\
        );

    \I__8910\ : InMux
    port map (
            O => \N__40489\,
            I => \N__40483\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__40486\,
            I => \N__40480\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__40483\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8907\ : Odrv4
    port map (
            O => \N__40480\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8906\ : InMux
    port map (
            O => \N__40475\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__8905\ : InMux
    port map (
            O => \N__40472\,
            I => \N__40468\
        );

    \I__8904\ : InMux
    port map (
            O => \N__40471\,
            I => \N__40465\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__40468\,
            I => \N__40462\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__40465\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8901\ : Odrv4
    port map (
            O => \N__40462\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8900\ : InMux
    port map (
            O => \N__40457\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__8899\ : InMux
    port map (
            O => \N__40454\,
            I => \N__40450\
        );

    \I__8898\ : InMux
    port map (
            O => \N__40453\,
            I => \N__40447\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__40450\,
            I => \N__40444\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__40447\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8895\ : Odrv4
    port map (
            O => \N__40444\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8894\ : InMux
    port map (
            O => \N__40439\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__8893\ : InMux
    port map (
            O => \N__40436\,
            I => \N__40433\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__40433\,
            I => \N__40430\
        );

    \I__8891\ : Span4Mux_h
    port map (
            O => \N__40430\,
            I => \N__40427\
        );

    \I__8890\ : Odrv4
    port map (
            O => \N__40427\,
            I => \phase_controller_inst2.stoper_tr.un6_running_12\
        );

    \I__8889\ : CascadeMux
    port map (
            O => \N__40424\,
            I => \N__40421\
        );

    \I__8888\ : InMux
    port map (
            O => \N__40421\,
            I => \N__40418\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__40418\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__8886\ : InMux
    port map (
            O => \N__40415\,
            I => \N__40412\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__40412\,
            I => \N__40409\
        );

    \I__8884\ : Span4Mux_h
    port map (
            O => \N__40409\,
            I => \N__40406\
        );

    \I__8883\ : Odrv4
    port map (
            O => \N__40406\,
            I => \phase_controller_inst2.stoper_tr.un6_running_13\
        );

    \I__8882\ : CascadeMux
    port map (
            O => \N__40403\,
            I => \N__40400\
        );

    \I__8881\ : InMux
    port map (
            O => \N__40400\,
            I => \N__40397\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__40397\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__8879\ : InMux
    port map (
            O => \N__40394\,
            I => \N__40391\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__40391\,
            I => \N__40388\
        );

    \I__8877\ : Span4Mux_h
    port map (
            O => \N__40388\,
            I => \N__40385\
        );

    \I__8876\ : Odrv4
    port map (
            O => \N__40385\,
            I => \phase_controller_inst2.stoper_tr.un6_running_14\
        );

    \I__8875\ : CascadeMux
    port map (
            O => \N__40382\,
            I => \N__40379\
        );

    \I__8874\ : InMux
    port map (
            O => \N__40379\,
            I => \N__40376\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__40376\,
            I => \N__40373\
        );

    \I__8872\ : Odrv4
    port map (
            O => \N__40373\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__8871\ : InMux
    port map (
            O => \N__40370\,
            I => \N__40367\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__40367\,
            I => \N__40364\
        );

    \I__8869\ : Span4Mux_v
    port map (
            O => \N__40364\,
            I => \N__40361\
        );

    \I__8868\ : Odrv4
    port map (
            O => \N__40361\,
            I => \phase_controller_inst2.stoper_tr.un6_running_15\
        );

    \I__8867\ : CascadeMux
    port map (
            O => \N__40358\,
            I => \N__40355\
        );

    \I__8866\ : InMux
    port map (
            O => \N__40355\,
            I => \N__40352\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__40352\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__8864\ : InMux
    port map (
            O => \N__40349\,
            I => \N__40346\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__40346\,
            I => \N__40343\
        );

    \I__8862\ : Span12Mux_h
    port map (
            O => \N__40343\,
            I => \N__40340\
        );

    \I__8861\ : Odrv12
    port map (
            O => \N__40340\,
            I => \phase_controller_inst2.stoper_tr.un6_running_16\
        );

    \I__8860\ : CascadeMux
    port map (
            O => \N__40337\,
            I => \N__40334\
        );

    \I__8859\ : InMux
    port map (
            O => \N__40334\,
            I => \N__40331\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__40331\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\
        );

    \I__8857\ : InMux
    port map (
            O => \N__40328\,
            I => \N__40325\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__40325\,
            I => \N__40322\
        );

    \I__8855\ : Span4Mux_h
    port map (
            O => \N__40322\,
            I => \N__40319\
        );

    \I__8854\ : Odrv4
    port map (
            O => \N__40319\,
            I => \phase_controller_inst2.stoper_tr.un6_running_17\
        );

    \I__8853\ : CascadeMux
    port map (
            O => \N__40316\,
            I => \N__40313\
        );

    \I__8852\ : InMux
    port map (
            O => \N__40313\,
            I => \N__40310\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__40310\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\
        );

    \I__8850\ : InMux
    port map (
            O => \N__40307\,
            I => \N__40304\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__40304\,
            I => \N__40301\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__40301\,
            I => \N__40298\
        );

    \I__8847\ : Odrv4
    port map (
            O => \N__40298\,
            I => \phase_controller_inst2.stoper_tr.un6_running_18\
        );

    \I__8846\ : CascadeMux
    port map (
            O => \N__40295\,
            I => \N__40292\
        );

    \I__8845\ : InMux
    port map (
            O => \N__40292\,
            I => \N__40289\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__40289\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\
        );

    \I__8843\ : InMux
    port map (
            O => \N__40286\,
            I => \N__40283\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__40283\,
            I => \N__40280\
        );

    \I__8841\ : Span4Mux_v
    port map (
            O => \N__40280\,
            I => \N__40277\
        );

    \I__8840\ : Odrv4
    port map (
            O => \N__40277\,
            I => \phase_controller_inst2.stoper_tr.un6_running_19\
        );

    \I__8839\ : CascadeMux
    port map (
            O => \N__40274\,
            I => \N__40271\
        );

    \I__8838\ : InMux
    port map (
            O => \N__40271\,
            I => \N__40268\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__40268\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\
        );

    \I__8836\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40262\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__40262\,
            I => \N__40259\
        );

    \I__8834\ : Span4Mux_v
    port map (
            O => \N__40259\,
            I => \N__40256\
        );

    \I__8833\ : Odrv4
    port map (
            O => \N__40256\,
            I => \phase_controller_inst2.stoper_tr.un6_running_4\
        );

    \I__8832\ : CascadeMux
    port map (
            O => \N__40253\,
            I => \N__40250\
        );

    \I__8831\ : InMux
    port map (
            O => \N__40250\,
            I => \N__40247\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__40247\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__8829\ : InMux
    port map (
            O => \N__40244\,
            I => \N__40241\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__40241\,
            I => \N__40238\
        );

    \I__8827\ : Span4Mux_v
    port map (
            O => \N__40238\,
            I => \N__40235\
        );

    \I__8826\ : Odrv4
    port map (
            O => \N__40235\,
            I => \phase_controller_inst2.stoper_tr.un6_running_5\
        );

    \I__8825\ : CascadeMux
    port map (
            O => \N__40232\,
            I => \N__40229\
        );

    \I__8824\ : InMux
    port map (
            O => \N__40229\,
            I => \N__40226\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__40226\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__8822\ : InMux
    port map (
            O => \N__40223\,
            I => \N__40220\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40220\,
            I => \N__40217\
        );

    \I__8820\ : Span4Mux_h
    port map (
            O => \N__40217\,
            I => \N__40214\
        );

    \I__8819\ : Odrv4
    port map (
            O => \N__40214\,
            I => \phase_controller_inst2.stoper_tr.un6_running_6\
        );

    \I__8818\ : CascadeMux
    port map (
            O => \N__40211\,
            I => \N__40208\
        );

    \I__8817\ : InMux
    port map (
            O => \N__40208\,
            I => \N__40205\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__40205\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__8815\ : InMux
    port map (
            O => \N__40202\,
            I => \N__40199\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__40199\,
            I => \N__40196\
        );

    \I__8813\ : Span4Mux_v
    port map (
            O => \N__40196\,
            I => \N__40193\
        );

    \I__8812\ : Odrv4
    port map (
            O => \N__40193\,
            I => \phase_controller_inst2.stoper_tr.un6_running_7\
        );

    \I__8811\ : CascadeMux
    port map (
            O => \N__40190\,
            I => \N__40187\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40187\,
            I => \N__40184\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__40184\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__8808\ : InMux
    port map (
            O => \N__40181\,
            I => \N__40178\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__40178\,
            I => \N__40175\
        );

    \I__8806\ : Span4Mux_h
    port map (
            O => \N__40175\,
            I => \N__40172\
        );

    \I__8805\ : Odrv4
    port map (
            O => \N__40172\,
            I => \phase_controller_inst2.stoper_tr.un6_running_8\
        );

    \I__8804\ : CascadeMux
    port map (
            O => \N__40169\,
            I => \N__40166\
        );

    \I__8803\ : InMux
    port map (
            O => \N__40166\,
            I => \N__40163\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__40163\,
            I => \N__40160\
        );

    \I__8801\ : Odrv4
    port map (
            O => \N__40160\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__8800\ : InMux
    port map (
            O => \N__40157\,
            I => \N__40154\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__40154\,
            I => \N__40151\
        );

    \I__8798\ : Span4Mux_h
    port map (
            O => \N__40151\,
            I => \N__40148\
        );

    \I__8797\ : Odrv4
    port map (
            O => \N__40148\,
            I => \phase_controller_inst2.stoper_tr.un6_running_9\
        );

    \I__8796\ : CascadeMux
    port map (
            O => \N__40145\,
            I => \N__40142\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40142\,
            I => \N__40139\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40139\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__8793\ : InMux
    port map (
            O => \N__40136\,
            I => \N__40133\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__40133\,
            I => \N__40130\
        );

    \I__8791\ : Span4Mux_h
    port map (
            O => \N__40130\,
            I => \N__40127\
        );

    \I__8790\ : Odrv4
    port map (
            O => \N__40127\,
            I => \phase_controller_inst2.stoper_tr.un6_running_10\
        );

    \I__8789\ : CascadeMux
    port map (
            O => \N__40124\,
            I => \N__40121\
        );

    \I__8788\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40118\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__40118\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__8786\ : InMux
    port map (
            O => \N__40115\,
            I => \N__40112\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__40112\,
            I => \N__40109\
        );

    \I__8784\ : Span4Mux_h
    port map (
            O => \N__40109\,
            I => \N__40106\
        );

    \I__8783\ : Odrv4
    port map (
            O => \N__40106\,
            I => \phase_controller_inst2.stoper_tr.un6_running_11\
        );

    \I__8782\ : CascadeMux
    port map (
            O => \N__40103\,
            I => \N__40100\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40100\,
            I => \N__40097\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__40097\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__8779\ : CascadeMux
    port map (
            O => \N__40094\,
            I => \elapsed_time_ns_1_RNI3JIF91_0_29_cascade_\
        );

    \I__8778\ : InMux
    port map (
            O => \N__40091\,
            I => \N__40088\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__40088\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\
        );

    \I__8776\ : CascadeMux
    port map (
            O => \N__40085\,
            I => \N__40082\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40082\,
            I => \N__40077\
        );

    \I__8774\ : InMux
    port map (
            O => \N__40081\,
            I => \N__40070\
        );

    \I__8773\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40070\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__40077\,
            I => \N__40067\
        );

    \I__8771\ : InMux
    port map (
            O => \N__40076\,
            I => \N__40062\
        );

    \I__8770\ : InMux
    port map (
            O => \N__40075\,
            I => \N__40062\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__40070\,
            I => \N__40059\
        );

    \I__8768\ : Odrv4
    port map (
            O => \N__40067\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__40062\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__8766\ : Odrv4
    port map (
            O => \N__40059\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40052\,
            I => \N__40049\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__40049\,
            I => \N__40046\
        );

    \I__8763\ : Span4Mux_h
    port map (
            O => \N__40046\,
            I => \N__40043\
        );

    \I__8762\ : Odrv4
    port map (
            O => \N__40043\,
            I => \phase_controller_inst1.stoper_tr.un6_running_14\
        );

    \I__8761\ : InMux
    port map (
            O => \N__40040\,
            I => \N__40036\
        );

    \I__8760\ : InMux
    port map (
            O => \N__40039\,
            I => \N__40033\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__40036\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__40033\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__8757\ : CascadeMux
    port map (
            O => \N__40028\,
            I => \N__40025\
        );

    \I__8756\ : InMux
    port map (
            O => \N__40025\,
            I => \N__40021\
        );

    \I__8755\ : InMux
    port map (
            O => \N__40024\,
            I => \N__40018\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__40021\,
            I => \N__40014\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__40018\,
            I => \N__40011\
        );

    \I__8752\ : InMux
    port map (
            O => \N__40017\,
            I => \N__40008\
        );

    \I__8751\ : Odrv4
    port map (
            O => \N__40014\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__8750\ : Odrv4
    port map (
            O => \N__40011\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__40008\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__8748\ : CascadeMux
    port map (
            O => \N__40001\,
            I => \N__39994\
        );

    \I__8747\ : CascadeMux
    port map (
            O => \N__40000\,
            I => \N__39985\
        );

    \I__8746\ : CascadeMux
    port map (
            O => \N__39999\,
            I => \N__39982\
        );

    \I__8745\ : InMux
    port map (
            O => \N__39998\,
            I => \N__39977\
        );

    \I__8744\ : InMux
    port map (
            O => \N__39997\,
            I => \N__39977\
        );

    \I__8743\ : InMux
    port map (
            O => \N__39994\,
            I => \N__39974\
        );

    \I__8742\ : InMux
    port map (
            O => \N__39993\,
            I => \N__39971\
        );

    \I__8741\ : InMux
    port map (
            O => \N__39992\,
            I => \N__39964\
        );

    \I__8740\ : InMux
    port map (
            O => \N__39991\,
            I => \N__39964\
        );

    \I__8739\ : InMux
    port map (
            O => \N__39990\,
            I => \N__39964\
        );

    \I__8738\ : InMux
    port map (
            O => \N__39989\,
            I => \N__39955\
        );

    \I__8737\ : InMux
    port map (
            O => \N__39988\,
            I => \N__39955\
        );

    \I__8736\ : InMux
    port map (
            O => \N__39985\,
            I => \N__39955\
        );

    \I__8735\ : InMux
    port map (
            O => \N__39982\,
            I => \N__39955\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__39977\,
            I => \N__39950\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__39974\,
            I => \N__39950\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__39971\,
            I => \phase_controller_inst1.stoper_tr.N_241\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__39964\,
            I => \phase_controller_inst1.stoper_tr.N_241\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__39955\,
            I => \phase_controller_inst1.stoper_tr.N_241\
        );

    \I__8729\ : Odrv12
    port map (
            O => \N__39950\,
            I => \phase_controller_inst1.stoper_tr.N_241\
        );

    \I__8728\ : CascadeMux
    port map (
            O => \N__39941\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\
        );

    \I__8727\ : InMux
    port map (
            O => \N__39938\,
            I => \N__39935\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__39935\,
            I => \N__39932\
        );

    \I__8725\ : Span4Mux_h
    port map (
            O => \N__39932\,
            I => \N__39929\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__39929\,
            I => \phase_controller_inst1.stoper_tr.un6_running_13\
        );

    \I__8723\ : InMux
    port map (
            O => \N__39926\,
            I => \N__39923\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__39923\,
            I => \N__39920\
        );

    \I__8721\ : Span4Mux_h
    port map (
            O => \N__39920\,
            I => \N__39914\
        );

    \I__8720\ : InMux
    port map (
            O => \N__39919\,
            I => \N__39911\
        );

    \I__8719\ : InMux
    port map (
            O => \N__39918\,
            I => \N__39906\
        );

    \I__8718\ : InMux
    port map (
            O => \N__39917\,
            I => \N__39906\
        );

    \I__8717\ : Odrv4
    port map (
            O => \N__39914\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__39911\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__39906\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19\
        );

    \I__8714\ : InMux
    port map (
            O => \N__39899\,
            I => \N__39866\
        );

    \I__8713\ : InMux
    port map (
            O => \N__39898\,
            I => \N__39866\
        );

    \I__8712\ : InMux
    port map (
            O => \N__39897\,
            I => \N__39866\
        );

    \I__8711\ : InMux
    port map (
            O => \N__39896\,
            I => \N__39853\
        );

    \I__8710\ : InMux
    port map (
            O => \N__39895\,
            I => \N__39853\
        );

    \I__8709\ : InMux
    port map (
            O => \N__39894\,
            I => \N__39844\
        );

    \I__8708\ : InMux
    port map (
            O => \N__39893\,
            I => \N__39844\
        );

    \I__8707\ : InMux
    port map (
            O => \N__39892\,
            I => \N__39844\
        );

    \I__8706\ : InMux
    port map (
            O => \N__39891\,
            I => \N__39844\
        );

    \I__8705\ : InMux
    port map (
            O => \N__39890\,
            I => \N__39841\
        );

    \I__8704\ : InMux
    port map (
            O => \N__39889\,
            I => \N__39836\
        );

    \I__8703\ : InMux
    port map (
            O => \N__39888\,
            I => \N__39836\
        );

    \I__8702\ : InMux
    port map (
            O => \N__39887\,
            I => \N__39829\
        );

    \I__8701\ : InMux
    port map (
            O => \N__39886\,
            I => \N__39829\
        );

    \I__8700\ : InMux
    port map (
            O => \N__39885\,
            I => \N__39829\
        );

    \I__8699\ : InMux
    port map (
            O => \N__39884\,
            I => \N__39822\
        );

    \I__8698\ : InMux
    port map (
            O => \N__39883\,
            I => \N__39822\
        );

    \I__8697\ : InMux
    port map (
            O => \N__39882\,
            I => \N__39822\
        );

    \I__8696\ : InMux
    port map (
            O => \N__39881\,
            I => \N__39807\
        );

    \I__8695\ : InMux
    port map (
            O => \N__39880\,
            I => \N__39807\
        );

    \I__8694\ : InMux
    port map (
            O => \N__39879\,
            I => \N__39807\
        );

    \I__8693\ : InMux
    port map (
            O => \N__39878\,
            I => \N__39807\
        );

    \I__8692\ : InMux
    port map (
            O => \N__39877\,
            I => \N__39807\
        );

    \I__8691\ : InMux
    port map (
            O => \N__39876\,
            I => \N__39807\
        );

    \I__8690\ : InMux
    port map (
            O => \N__39875\,
            I => \N__39807\
        );

    \I__8689\ : InMux
    port map (
            O => \N__39874\,
            I => \N__39802\
        );

    \I__8688\ : InMux
    port map (
            O => \N__39873\,
            I => \N__39802\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__39866\,
            I => \N__39799\
        );

    \I__8686\ : InMux
    port map (
            O => \N__39865\,
            I => \N__39788\
        );

    \I__8685\ : InMux
    port map (
            O => \N__39864\,
            I => \N__39788\
        );

    \I__8684\ : InMux
    port map (
            O => \N__39863\,
            I => \N__39788\
        );

    \I__8683\ : InMux
    port map (
            O => \N__39862\,
            I => \N__39788\
        );

    \I__8682\ : InMux
    port map (
            O => \N__39861\,
            I => \N__39788\
        );

    \I__8681\ : InMux
    port map (
            O => \N__39860\,
            I => \N__39781\
        );

    \I__8680\ : InMux
    port map (
            O => \N__39859\,
            I => \N__39781\
        );

    \I__8679\ : InMux
    port map (
            O => \N__39858\,
            I => \N__39781\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__39853\,
            I => \N__39772\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__39844\,
            I => \N__39772\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__39841\,
            I => \N__39772\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__39836\,
            I => \N__39772\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__39829\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__39822\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__39807\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__39802\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__8670\ : Odrv4
    port map (
            O => \N__39799\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__39788\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__39781\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__8667\ : Odrv4
    port map (
            O => \N__39772\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__8666\ : CascadeMux
    port map (
            O => \N__39755\,
            I => \N__39748\
        );

    \I__8665\ : CascadeMux
    port map (
            O => \N__39754\,
            I => \N__39745\
        );

    \I__8664\ : InMux
    port map (
            O => \N__39753\,
            I => \N__39717\
        );

    \I__8663\ : InMux
    port map (
            O => \N__39752\,
            I => \N__39717\
        );

    \I__8662\ : InMux
    port map (
            O => \N__39751\,
            I => \N__39717\
        );

    \I__8661\ : InMux
    port map (
            O => \N__39748\,
            I => \N__39717\
        );

    \I__8660\ : InMux
    port map (
            O => \N__39745\,
            I => \N__39717\
        );

    \I__8659\ : InMux
    port map (
            O => \N__39744\,
            I => \N__39703\
        );

    \I__8658\ : InMux
    port map (
            O => \N__39743\,
            I => \N__39703\
        );

    \I__8657\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39703\
        );

    \I__8656\ : InMux
    port map (
            O => \N__39741\,
            I => \N__39703\
        );

    \I__8655\ : InMux
    port map (
            O => \N__39740\,
            I => \N__39703\
        );

    \I__8654\ : InMux
    port map (
            O => \N__39739\,
            I => \N__39698\
        );

    \I__8653\ : InMux
    port map (
            O => \N__39738\,
            I => \N__39698\
        );

    \I__8652\ : InMux
    port map (
            O => \N__39737\,
            I => \N__39691\
        );

    \I__8651\ : InMux
    port map (
            O => \N__39736\,
            I => \N__39691\
        );

    \I__8650\ : InMux
    port map (
            O => \N__39735\,
            I => \N__39691\
        );

    \I__8649\ : InMux
    port map (
            O => \N__39734\,
            I => \N__39688\
        );

    \I__8648\ : InMux
    port map (
            O => \N__39733\,
            I => \N__39685\
        );

    \I__8647\ : InMux
    port map (
            O => \N__39732\,
            I => \N__39678\
        );

    \I__8646\ : InMux
    port map (
            O => \N__39731\,
            I => \N__39678\
        );

    \I__8645\ : InMux
    port map (
            O => \N__39730\,
            I => \N__39678\
        );

    \I__8644\ : CascadeMux
    port map (
            O => \N__39729\,
            I => \N__39674\
        );

    \I__8643\ : CascadeMux
    port map (
            O => \N__39728\,
            I => \N__39670\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__39717\,
            I => \N__39667\
        );

    \I__8641\ : InMux
    port map (
            O => \N__39716\,
            I => \N__39660\
        );

    \I__8640\ : InMux
    port map (
            O => \N__39715\,
            I => \N__39660\
        );

    \I__8639\ : InMux
    port map (
            O => \N__39714\,
            I => \N__39660\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__39703\,
            I => \N__39653\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__39698\,
            I => \N__39653\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__39691\,
            I => \N__39653\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__39688\,
            I => \N__39646\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__39685\,
            I => \N__39646\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__39678\,
            I => \N__39646\
        );

    \I__8632\ : InMux
    port map (
            O => \N__39677\,
            I => \N__39643\
        );

    \I__8631\ : InMux
    port map (
            O => \N__39674\,
            I => \N__39636\
        );

    \I__8630\ : InMux
    port map (
            O => \N__39673\,
            I => \N__39636\
        );

    \I__8629\ : InMux
    port map (
            O => \N__39670\,
            I => \N__39636\
        );

    \I__8628\ : Span4Mux_v
    port map (
            O => \N__39667\,
            I => \N__39633\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__39660\,
            I => \N__39628\
        );

    \I__8626\ : Span4Mux_h
    port map (
            O => \N__39653\,
            I => \N__39628\
        );

    \I__8625\ : Span4Mux_v
    port map (
            O => \N__39646\,
            I => \N__39623\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__39643\,
            I => \N__39623\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__39636\,
            I => \N__39620\
        );

    \I__8622\ : Odrv4
    port map (
            O => \N__39633\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8621\ : Odrv4
    port map (
            O => \N__39628\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8620\ : Odrv4
    port map (
            O => \N__39623\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8619\ : Odrv12
    port map (
            O => \N__39620\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8618\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39608\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__39608\,
            I => \N__39605\
        );

    \I__8616\ : Span4Mux_h
    port map (
            O => \N__39605\,
            I => \N__39602\
        );

    \I__8615\ : Odrv4
    port map (
            O => \N__39602\,
            I => \phase_controller_inst1.stoper_tr.un6_running_19\
        );

    \I__8614\ : CEMux
    port map (
            O => \N__39599\,
            I => \N__39594\
        );

    \I__8613\ : CEMux
    port map (
            O => \N__39598\,
            I => \N__39591\
        );

    \I__8612\ : CEMux
    port map (
            O => \N__39597\,
            I => \N__39582\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__39594\,
            I => \N__39575\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__39591\,
            I => \N__39572\
        );

    \I__8609\ : InMux
    port map (
            O => \N__39590\,
            I => \N__39563\
        );

    \I__8608\ : InMux
    port map (
            O => \N__39589\,
            I => \N__39563\
        );

    \I__8607\ : InMux
    port map (
            O => \N__39588\,
            I => \N__39563\
        );

    \I__8606\ : InMux
    port map (
            O => \N__39587\,
            I => \N__39563\
        );

    \I__8605\ : InMux
    port map (
            O => \N__39586\,
            I => \N__39560\
        );

    \I__8604\ : CEMux
    port map (
            O => \N__39585\,
            I => \N__39557\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__39582\,
            I => \N__39554\
        );

    \I__8602\ : InMux
    port map (
            O => \N__39581\,
            I => \N__39535\
        );

    \I__8601\ : InMux
    port map (
            O => \N__39580\,
            I => \N__39535\
        );

    \I__8600\ : InMux
    port map (
            O => \N__39579\,
            I => \N__39535\
        );

    \I__8599\ : InMux
    port map (
            O => \N__39578\,
            I => \N__39535\
        );

    \I__8598\ : Span4Mux_v
    port map (
            O => \N__39575\,
            I => \N__39532\
        );

    \I__8597\ : Span4Mux_h
    port map (
            O => \N__39572\,
            I => \N__39529\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__39563\,
            I => \N__39524\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__39560\,
            I => \N__39524\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__39557\,
            I => \N__39519\
        );

    \I__8593\ : Span4Mux_h
    port map (
            O => \N__39554\,
            I => \N__39519\
        );

    \I__8592\ : InMux
    port map (
            O => \N__39553\,
            I => \N__39512\
        );

    \I__8591\ : InMux
    port map (
            O => \N__39552\,
            I => \N__39512\
        );

    \I__8590\ : InMux
    port map (
            O => \N__39551\,
            I => \N__39512\
        );

    \I__8589\ : InMux
    port map (
            O => \N__39550\,
            I => \N__39509\
        );

    \I__8588\ : InMux
    port map (
            O => \N__39549\,
            I => \N__39504\
        );

    \I__8587\ : InMux
    port map (
            O => \N__39548\,
            I => \N__39504\
        );

    \I__8586\ : InMux
    port map (
            O => \N__39547\,
            I => \N__39495\
        );

    \I__8585\ : InMux
    port map (
            O => \N__39546\,
            I => \N__39495\
        );

    \I__8584\ : InMux
    port map (
            O => \N__39545\,
            I => \N__39495\
        );

    \I__8583\ : InMux
    port map (
            O => \N__39544\,
            I => \N__39495\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__39535\,
            I => \N__39490\
        );

    \I__8581\ : Span4Mux_h
    port map (
            O => \N__39532\,
            I => \N__39490\
        );

    \I__8580\ : Span4Mux_v
    port map (
            O => \N__39529\,
            I => \N__39485\
        );

    \I__8579\ : Span4Mux_h
    port map (
            O => \N__39524\,
            I => \N__39485\
        );

    \I__8578\ : Span4Mux_h
    port map (
            O => \N__39519\,
            I => \N__39482\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__39512\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__39509\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__39504\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__39495\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__8573\ : Odrv4
    port map (
            O => \N__39490\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__8572\ : Odrv4
    port map (
            O => \N__39485\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__8571\ : Odrv4
    port map (
            O => \N__39482\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__8570\ : InMux
    port map (
            O => \N__39467\,
            I => \N__39464\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__39464\,
            I => \N__39461\
        );

    \I__8568\ : Span4Mux_h
    port map (
            O => \N__39461\,
            I => \N__39458\
        );

    \I__8567\ : Odrv4
    port map (
            O => \N__39458\,
            I => \phase_controller_inst2.stoper_tr.un6_running_1\
        );

    \I__8566\ : CascadeMux
    port map (
            O => \N__39455\,
            I => \N__39452\
        );

    \I__8565\ : InMux
    port map (
            O => \N__39452\,
            I => \N__39449\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__39449\,
            I => \N__39446\
        );

    \I__8563\ : Odrv4
    port map (
            O => \N__39446\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__8562\ : InMux
    port map (
            O => \N__39443\,
            I => \N__39440\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__39440\,
            I => \N__39437\
        );

    \I__8560\ : Span4Mux_h
    port map (
            O => \N__39437\,
            I => \N__39434\
        );

    \I__8559\ : Odrv4
    port map (
            O => \N__39434\,
            I => \phase_controller_inst2.stoper_tr.un6_running_2\
        );

    \I__8558\ : CascadeMux
    port map (
            O => \N__39431\,
            I => \N__39428\
        );

    \I__8557\ : InMux
    port map (
            O => \N__39428\,
            I => \N__39425\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__39425\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__8555\ : InMux
    port map (
            O => \N__39422\,
            I => \N__39419\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__39419\,
            I => \N__39416\
        );

    \I__8553\ : Span4Mux_v
    port map (
            O => \N__39416\,
            I => \N__39413\
        );

    \I__8552\ : Odrv4
    port map (
            O => \N__39413\,
            I => \phase_controller_inst2.stoper_tr.un6_running_3\
        );

    \I__8551\ : CascadeMux
    port map (
            O => \N__39410\,
            I => \N__39407\
        );

    \I__8550\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39404\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__39404\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__8548\ : CascadeMux
    port map (
            O => \N__39401\,
            I => \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\
        );

    \I__8547\ : InMux
    port map (
            O => \N__39398\,
            I => \N__39394\
        );

    \I__8546\ : InMux
    port map (
            O => \N__39397\,
            I => \N__39391\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__39394\,
            I => \elapsed_time_ns_1_RNIRAIF91_0_21\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__39391\,
            I => \elapsed_time_ns_1_RNIRAIF91_0_21\
        );

    \I__8543\ : CascadeMux
    port map (
            O => \N__39386\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_\
        );

    \I__8542\ : InMux
    port map (
            O => \N__39383\,
            I => \N__39379\
        );

    \I__8541\ : InMux
    port map (
            O => \N__39382\,
            I => \N__39376\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__39379\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__39376\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__8538\ : InMux
    port map (
            O => \N__39371\,
            I => \N__39367\
        );

    \I__8537\ : InMux
    port map (
            O => \N__39370\,
            I => \N__39364\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__39367\,
            I => \N__39360\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__39364\,
            I => \N__39357\
        );

    \I__8534\ : CascadeMux
    port map (
            O => \N__39363\,
            I => \N__39353\
        );

    \I__8533\ : Span4Mux_v
    port map (
            O => \N__39360\,
            I => \N__39348\
        );

    \I__8532\ : Span4Mux_v
    port map (
            O => \N__39357\,
            I => \N__39348\
        );

    \I__8531\ : InMux
    port map (
            O => \N__39356\,
            I => \N__39345\
        );

    \I__8530\ : InMux
    port map (
            O => \N__39353\,
            I => \N__39342\
        );

    \I__8529\ : Sp12to4
    port map (
            O => \N__39348\,
            I => \N__39337\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__39345\,
            I => \N__39337\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__39342\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__8526\ : Odrv12
    port map (
            O => \N__39337\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__8525\ : CascadeMux
    port map (
            O => \N__39332\,
            I => \N__39328\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39331\,
            I => \N__39325\
        );

    \I__8523\ : InMux
    port map (
            O => \N__39328\,
            I => \N__39322\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__39325\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__39322\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__8520\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39311\
        );

    \I__8519\ : InMux
    port map (
            O => \N__39316\,
            I => \N__39311\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__39311\,
            I => \delay_measurement_inst.delay_tr_timer.N_347\
        );

    \I__8517\ : InMux
    port map (
            O => \N__39308\,
            I => \N__39305\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__39305\,
            I => \N__39301\
        );

    \I__8515\ : InMux
    port map (
            O => \N__39304\,
            I => \N__39298\
        );

    \I__8514\ : Odrv4
    port map (
            O => \N__39301\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__39298\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__8512\ : CascadeMux
    port map (
            O => \N__39293\,
            I => \N__39290\
        );

    \I__8511\ : InMux
    port map (
            O => \N__39290\,
            I => \N__39287\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__39287\,
            I => \N__39283\
        );

    \I__8509\ : InMux
    port map (
            O => \N__39286\,
            I => \N__39280\
        );

    \I__8508\ : Odrv4
    port map (
            O => \N__39283\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__39280\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__8506\ : InMux
    port map (
            O => \N__39275\,
            I => \N__39269\
        );

    \I__8505\ : InMux
    port map (
            O => \N__39274\,
            I => \N__39269\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__39269\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__8503\ : CascadeMux
    port map (
            O => \N__39266\,
            I => \N__39263\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39263\,
            I => \N__39259\
        );

    \I__8501\ : InMux
    port map (
            O => \N__39262\,
            I => \N__39256\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__39259\,
            I => \N__39253\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__39256\,
            I => \N__39247\
        );

    \I__8498\ : Span4Mux_v
    port map (
            O => \N__39253\,
            I => \N__39247\
        );

    \I__8497\ : InMux
    port map (
            O => \N__39252\,
            I => \N__39244\
        );

    \I__8496\ : Odrv4
    port map (
            O => \N__39247\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__39244\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__8494\ : CascadeMux
    port map (
            O => \N__39239\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11_cascade_\
        );

    \I__8493\ : CascadeMux
    port map (
            O => \N__39236\,
            I => \N__39233\
        );

    \I__8492\ : InMux
    port map (
            O => \N__39233\,
            I => \N__39228\
        );

    \I__8491\ : InMux
    port map (
            O => \N__39232\,
            I => \N__39225\
        );

    \I__8490\ : CascadeMux
    port map (
            O => \N__39231\,
            I => \N__39222\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__39228\,
            I => \N__39217\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__39225\,
            I => \N__39217\
        );

    \I__8487\ : InMux
    port map (
            O => \N__39222\,
            I => \N__39213\
        );

    \I__8486\ : Span4Mux_v
    port map (
            O => \N__39217\,
            I => \N__39210\
        );

    \I__8485\ : InMux
    port map (
            O => \N__39216\,
            I => \N__39207\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__39213\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__8483\ : Odrv4
    port map (
            O => \N__39210\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__39207\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__8481\ : CascadeMux
    port map (
            O => \N__39200\,
            I => \N__39195\
        );

    \I__8480\ : InMux
    port map (
            O => \N__39199\,
            I => \N__39192\
        );

    \I__8479\ : InMux
    port map (
            O => \N__39198\,
            I => \N__39189\
        );

    \I__8478\ : InMux
    port map (
            O => \N__39195\,
            I => \N__39186\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__39192\,
            I => \N__39181\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39189\,
            I => \N__39181\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__39186\,
            I => \N__39178\
        );

    \I__8474\ : Span4Mux_v
    port map (
            O => \N__39181\,
            I => \N__39173\
        );

    \I__8473\ : Span4Mux_v
    port map (
            O => \N__39178\,
            I => \N__39173\
        );

    \I__8472\ : Odrv4
    port map (
            O => \N__39173\,
            I => \phase_controller_inst1.stoper_tr.N_244\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39170\,
            I => \N__39164\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39169\,
            I => \N__39164\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__39164\,
            I => \N__39161\
        );

    \I__8468\ : Odrv4
    port map (
            O => \N__39161\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39158\,
            I => \N__39155\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__39155\,
            I => \elapsed_time_ns_1_RNI3JIF91_0_29\
        );

    \I__8465\ : CascadeMux
    port map (
            O => \N__39152\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\
        );

    \I__8464\ : CascadeMux
    port map (
            O => \N__39149\,
            I => \delay_measurement_inst.delay_tr_timer.N_358_cascade_\
        );

    \I__8463\ : InMux
    port map (
            O => \N__39146\,
            I => \N__39143\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__39143\,
            I => \delay_measurement_inst.delay_tr_timer.N_381\
        );

    \I__8461\ : InMux
    port map (
            O => \N__39140\,
            I => \N__39130\
        );

    \I__8460\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39127\
        );

    \I__8459\ : InMux
    port map (
            O => \N__39138\,
            I => \N__39124\
        );

    \I__8458\ : InMux
    port map (
            O => \N__39137\,
            I => \N__39121\
        );

    \I__8457\ : InMux
    port map (
            O => \N__39136\,
            I => \N__39118\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39135\,
            I => \N__39113\
        );

    \I__8455\ : InMux
    port map (
            O => \N__39134\,
            I => \N__39113\
        );

    \I__8454\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39110\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__39130\,
            I => \N__39104\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__39127\,
            I => \N__39104\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__39124\,
            I => \N__39099\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__39121\,
            I => \N__39099\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__39118\,
            I => \N__39094\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39113\,
            I => \N__39094\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__39110\,
            I => \N__39091\
        );

    \I__8446\ : InMux
    port map (
            O => \N__39109\,
            I => \N__39088\
        );

    \I__8445\ : Span4Mux_h
    port map (
            O => \N__39104\,
            I => \N__39085\
        );

    \I__8444\ : Span4Mux_h
    port map (
            O => \N__39099\,
            I => \N__39082\
        );

    \I__8443\ : Span4Mux_h
    port map (
            O => \N__39094\,
            I => \N__39079\
        );

    \I__8442\ : Odrv12
    port map (
            O => \N__39091\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__39088\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__8440\ : Odrv4
    port map (
            O => \N__39085\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__8439\ : Odrv4
    port map (
            O => \N__39082\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__8438\ : Odrv4
    port map (
            O => \N__39079\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__8437\ : InMux
    port map (
            O => \N__39068\,
            I => \N__39065\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__39065\,
            I => \N__39059\
        );

    \I__8435\ : InMux
    port map (
            O => \N__39064\,
            I => \N__39056\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39063\,
            I => \N__39051\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39062\,
            I => \N__39051\
        );

    \I__8432\ : Odrv4
    port map (
            O => \N__39059\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__39056\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__39051\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__8429\ : InMux
    port map (
            O => \N__39044\,
            I => \N__39041\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__39041\,
            I => \N__39037\
        );

    \I__8427\ : CascadeMux
    port map (
            O => \N__39040\,
            I => \N__39034\
        );

    \I__8426\ : Span4Mux_v
    port map (
            O => \N__39037\,
            I => \N__39030\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39034\,
            I => \N__39025\
        );

    \I__8424\ : InMux
    port map (
            O => \N__39033\,
            I => \N__39025\
        );

    \I__8423\ : Odrv4
    port map (
            O => \N__39030\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__39025\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__8421\ : CascadeMux
    port map (
            O => \N__39020\,
            I => \delay_measurement_inst.delay_tr_timer.N_348_cascade_\
        );

    \I__8420\ : InMux
    port map (
            O => \N__39017\,
            I => \N__39014\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__39014\,
            I => \N__39008\
        );

    \I__8418\ : InMux
    port map (
            O => \N__39013\,
            I => \N__39005\
        );

    \I__8417\ : InMux
    port map (
            O => \N__39012\,
            I => \N__39000\
        );

    \I__8416\ : InMux
    port map (
            O => \N__39011\,
            I => \N__39000\
        );

    \I__8415\ : Odrv4
    port map (
            O => \N__39008\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__39005\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__39000\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__8412\ : InMux
    port map (
            O => \N__38993\,
            I => \N__38984\
        );

    \I__8411\ : InMux
    port map (
            O => \N__38992\,
            I => \N__38984\
        );

    \I__8410\ : InMux
    port map (
            O => \N__38991\,
            I => \N__38984\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__38984\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__8408\ : InMux
    port map (
            O => \N__38981\,
            I => \N__38978\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__38978\,
            I => \N__38973\
        );

    \I__8406\ : InMux
    port map (
            O => \N__38977\,
            I => \N__38970\
        );

    \I__8405\ : InMux
    port map (
            O => \N__38976\,
            I => \N__38967\
        );

    \I__8404\ : Span4Mux_h
    port map (
            O => \N__38973\,
            I => \N__38961\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__38970\,
            I => \N__38961\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__38967\,
            I => \N__38958\
        );

    \I__8401\ : InMux
    port map (
            O => \N__38966\,
            I => \N__38955\
        );

    \I__8400\ : Span4Mux_v
    port map (
            O => \N__38961\,
            I => \N__38952\
        );

    \I__8399\ : Span4Mux_v
    port map (
            O => \N__38958\,
            I => \N__38949\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__38955\,
            I => \N__38946\
        );

    \I__8397\ : Odrv4
    port map (
            O => \N__38952\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__8396\ : Odrv4
    port map (
            O => \N__38949\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__8395\ : Odrv12
    port map (
            O => \N__38946\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__8394\ : InMux
    port map (
            O => \N__38939\,
            I => \N__38936\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__38936\,
            I => \elapsed_time_ns_1_RNITCIF91_0_23\
        );

    \I__8392\ : CascadeMux
    port map (
            O => \N__38933\,
            I => \N__38930\
        );

    \I__8391\ : InMux
    port map (
            O => \N__38930\,
            I => \N__38926\
        );

    \I__8390\ : InMux
    port map (
            O => \N__38929\,
            I => \N__38923\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__38926\,
            I => \N__38920\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__38923\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__8387\ : Odrv4
    port map (
            O => \N__38920\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__8386\ : InMux
    port map (
            O => \N__38915\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__8385\ : InMux
    port map (
            O => \N__38912\,
            I => \N__38888\
        );

    \I__8384\ : InMux
    port map (
            O => \N__38911\,
            I => \N__38888\
        );

    \I__8383\ : InMux
    port map (
            O => \N__38910\,
            I => \N__38888\
        );

    \I__8382\ : InMux
    port map (
            O => \N__38909\,
            I => \N__38888\
        );

    \I__8381\ : InMux
    port map (
            O => \N__38908\,
            I => \N__38879\
        );

    \I__8380\ : InMux
    port map (
            O => \N__38907\,
            I => \N__38879\
        );

    \I__8379\ : InMux
    port map (
            O => \N__38906\,
            I => \N__38879\
        );

    \I__8378\ : InMux
    port map (
            O => \N__38905\,
            I => \N__38879\
        );

    \I__8377\ : InMux
    port map (
            O => \N__38904\,
            I => \N__38856\
        );

    \I__8376\ : InMux
    port map (
            O => \N__38903\,
            I => \N__38856\
        );

    \I__8375\ : InMux
    port map (
            O => \N__38902\,
            I => \N__38856\
        );

    \I__8374\ : InMux
    port map (
            O => \N__38901\,
            I => \N__38856\
        );

    \I__8373\ : InMux
    port map (
            O => \N__38900\,
            I => \N__38847\
        );

    \I__8372\ : InMux
    port map (
            O => \N__38899\,
            I => \N__38847\
        );

    \I__8371\ : InMux
    port map (
            O => \N__38898\,
            I => \N__38847\
        );

    \I__8370\ : InMux
    port map (
            O => \N__38897\,
            I => \N__38847\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__38888\,
            I => \N__38844\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__38879\,
            I => \N__38841\
        );

    \I__8367\ : InMux
    port map (
            O => \N__38878\,
            I => \N__38836\
        );

    \I__8366\ : InMux
    port map (
            O => \N__38877\,
            I => \N__38836\
        );

    \I__8365\ : InMux
    port map (
            O => \N__38876\,
            I => \N__38827\
        );

    \I__8364\ : InMux
    port map (
            O => \N__38875\,
            I => \N__38827\
        );

    \I__8363\ : InMux
    port map (
            O => \N__38874\,
            I => \N__38827\
        );

    \I__8362\ : InMux
    port map (
            O => \N__38873\,
            I => \N__38827\
        );

    \I__8361\ : InMux
    port map (
            O => \N__38872\,
            I => \N__38818\
        );

    \I__8360\ : InMux
    port map (
            O => \N__38871\,
            I => \N__38818\
        );

    \I__8359\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38818\
        );

    \I__8358\ : InMux
    port map (
            O => \N__38869\,
            I => \N__38818\
        );

    \I__8357\ : InMux
    port map (
            O => \N__38868\,
            I => \N__38809\
        );

    \I__8356\ : InMux
    port map (
            O => \N__38867\,
            I => \N__38809\
        );

    \I__8355\ : InMux
    port map (
            O => \N__38866\,
            I => \N__38809\
        );

    \I__8354\ : InMux
    port map (
            O => \N__38865\,
            I => \N__38809\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__38856\,
            I => \N__38804\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__38847\,
            I => \N__38804\
        );

    \I__8351\ : Span4Mux_h
    port map (
            O => \N__38844\,
            I => \N__38799\
        );

    \I__8350\ : Span4Mux_h
    port map (
            O => \N__38841\,
            I => \N__38799\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__38836\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__38827\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__38818\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__38809\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8345\ : Odrv4
    port map (
            O => \N__38804\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8344\ : Odrv4
    port map (
            O => \N__38799\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8343\ : InMux
    port map (
            O => \N__38786\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__8342\ : InMux
    port map (
            O => \N__38783\,
            I => \N__38779\
        );

    \I__8341\ : InMux
    port map (
            O => \N__38782\,
            I => \N__38776\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__38779\,
            I => \N__38773\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__38776\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__8338\ : Odrv4
    port map (
            O => \N__38773\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__8337\ : CEMux
    port map (
            O => \N__38768\,
            I => \N__38763\
        );

    \I__8336\ : CEMux
    port map (
            O => \N__38767\,
            I => \N__38760\
        );

    \I__8335\ : CEMux
    port map (
            O => \N__38766\,
            I => \N__38757\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__38763\,
            I => \N__38754\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__38760\,
            I => \N__38751\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__38757\,
            I => \N__38747\
        );

    \I__8331\ : Span4Mux_v
    port map (
            O => \N__38754\,
            I => \N__38742\
        );

    \I__8330\ : Span4Mux_h
    port map (
            O => \N__38751\,
            I => \N__38742\
        );

    \I__8329\ : CEMux
    port map (
            O => \N__38750\,
            I => \N__38739\
        );

    \I__8328\ : Span4Mux_v
    port map (
            O => \N__38747\,
            I => \N__38732\
        );

    \I__8327\ : Span4Mux_h
    port map (
            O => \N__38742\,
            I => \N__38732\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__38739\,
            I => \N__38732\
        );

    \I__8325\ : Span4Mux_v
    port map (
            O => \N__38732\,
            I => \N__38729\
        );

    \I__8324\ : Odrv4
    port map (
            O => \N__38729\,
            I => \current_shift_inst.timer_s1.N_167_i\
        );

    \I__8323\ : CascadeMux
    port map (
            O => \N__38726\,
            I => \N__38722\
        );

    \I__8322\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38719\
        );

    \I__8321\ : InMux
    port map (
            O => \N__38722\,
            I => \N__38716\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__38719\,
            I => \N__38710\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__38716\,
            I => \N__38710\
        );

    \I__8318\ : InMux
    port map (
            O => \N__38715\,
            I => \N__38707\
        );

    \I__8317\ : Span4Mux_v
    port map (
            O => \N__38710\,
            I => \N__38704\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__38707\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8315\ : Odrv4
    port map (
            O => \N__38704\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8314\ : CEMux
    port map (
            O => \N__38699\,
            I => \N__38681\
        );

    \I__8313\ : CEMux
    port map (
            O => \N__38698\,
            I => \N__38681\
        );

    \I__8312\ : CEMux
    port map (
            O => \N__38697\,
            I => \N__38681\
        );

    \I__8311\ : CEMux
    port map (
            O => \N__38696\,
            I => \N__38681\
        );

    \I__8310\ : CEMux
    port map (
            O => \N__38695\,
            I => \N__38681\
        );

    \I__8309\ : CEMux
    port map (
            O => \N__38694\,
            I => \N__38681\
        );

    \I__8308\ : GlobalMux
    port map (
            O => \N__38681\,
            I => \N__38678\
        );

    \I__8307\ : gio2CtrlBuf
    port map (
            O => \N__38678\,
            I => \delay_measurement_inst.delay_tr_timer.N_434_i_g\
        );

    \I__8306\ : CascadeMux
    port map (
            O => \N__38675\,
            I => \N__38671\
        );

    \I__8305\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38665\
        );

    \I__8304\ : InMux
    port map (
            O => \N__38671\,
            I => \N__38665\
        );

    \I__8303\ : InMux
    port map (
            O => \N__38670\,
            I => \N__38662\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__38665\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__38662\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__8300\ : InMux
    port map (
            O => \N__38657\,
            I => \N__38654\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__38654\,
            I => \N__38650\
        );

    \I__8298\ : CascadeMux
    port map (
            O => \N__38653\,
            I => \N__38647\
        );

    \I__8297\ : Span4Mux_h
    port map (
            O => \N__38650\,
            I => \N__38644\
        );

    \I__8296\ : InMux
    port map (
            O => \N__38647\,
            I => \N__38641\
        );

    \I__8295\ : Odrv4
    port map (
            O => \N__38644\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__38641\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__8293\ : InMux
    port map (
            O => \N__38636\,
            I => \N__38632\
        );

    \I__8292\ : InMux
    port map (
            O => \N__38635\,
            I => \N__38629\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__38632\,
            I => \delay_measurement_inst.delay_tr_timer.N_341\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__38629\,
            I => \delay_measurement_inst.delay_tr_timer.N_341\
        );

    \I__8289\ : CascadeMux
    port map (
            O => \N__38624\,
            I => \N__38620\
        );

    \I__8288\ : InMux
    port map (
            O => \N__38623\,
            I => \N__38616\
        );

    \I__8287\ : InMux
    port map (
            O => \N__38620\,
            I => \N__38611\
        );

    \I__8286\ : InMux
    port map (
            O => \N__38619\,
            I => \N__38611\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__38616\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__38611\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__8283\ : CascadeMux
    port map (
            O => \N__38606\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\
        );

    \I__8282\ : InMux
    port map (
            O => \N__38603\,
            I => \N__38600\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__38600\,
            I => \N__38596\
        );

    \I__8280\ : InMux
    port map (
            O => \N__38599\,
            I => \N__38593\
        );

    \I__8279\ : Span4Mux_v
    port map (
            O => \N__38596\,
            I => \N__38585\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__38593\,
            I => \N__38585\
        );

    \I__8277\ : InMux
    port map (
            O => \N__38592\,
            I => \N__38580\
        );

    \I__8276\ : InMux
    port map (
            O => \N__38591\,
            I => \N__38580\
        );

    \I__8275\ : InMux
    port map (
            O => \N__38590\,
            I => \N__38577\
        );

    \I__8274\ : Span4Mux_h
    port map (
            O => \N__38585\,
            I => \N__38574\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__38580\,
            I => \N__38571\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__38577\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__8271\ : Odrv4
    port map (
            O => \N__38574\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__8270\ : Odrv12
    port map (
            O => \N__38571\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__8269\ : CascadeMux
    port map (
            O => \N__38564\,
            I => \delay_measurement_inst.delay_tr_timer.N_381_cascade_\
        );

    \I__8268\ : InMux
    port map (
            O => \N__38561\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__8267\ : CascadeMux
    port map (
            O => \N__38558\,
            I => \N__38554\
        );

    \I__8266\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38550\
        );

    \I__8265\ : InMux
    port map (
            O => \N__38554\,
            I => \N__38547\
        );

    \I__8264\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38544\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__38550\,
            I => \N__38539\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__38547\,
            I => \N__38539\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__38544\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__8260\ : Odrv4
    port map (
            O => \N__38539\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__8259\ : InMux
    port map (
            O => \N__38534\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__8258\ : CascadeMux
    port map (
            O => \N__38531\,
            I => \N__38528\
        );

    \I__8257\ : InMux
    port map (
            O => \N__38528\,
            I => \N__38523\
        );

    \I__8256\ : InMux
    port map (
            O => \N__38527\,
            I => \N__38520\
        );

    \I__8255\ : InMux
    port map (
            O => \N__38526\,
            I => \N__38517\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__38523\,
            I => \N__38512\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__38520\,
            I => \N__38512\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__38517\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__8251\ : Odrv4
    port map (
            O => \N__38512\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__8250\ : InMux
    port map (
            O => \N__38507\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__8249\ : CascadeMux
    port map (
            O => \N__38504\,
            I => \N__38500\
        );

    \I__8248\ : CascadeMux
    port map (
            O => \N__38503\,
            I => \N__38497\
        );

    \I__8247\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38491\
        );

    \I__8246\ : InMux
    port map (
            O => \N__38497\,
            I => \N__38491\
        );

    \I__8245\ : InMux
    port map (
            O => \N__38496\,
            I => \N__38488\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__38491\,
            I => \N__38485\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__38488\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__8242\ : Odrv4
    port map (
            O => \N__38485\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__8241\ : InMux
    port map (
            O => \N__38480\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__8240\ : InMux
    port map (
            O => \N__38477\,
            I => \N__38470\
        );

    \I__8239\ : InMux
    port map (
            O => \N__38476\,
            I => \N__38470\
        );

    \I__8238\ : InMux
    port map (
            O => \N__38475\,
            I => \N__38467\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__38470\,
            I => \N__38464\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__38467\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__8235\ : Odrv4
    port map (
            O => \N__38464\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__8234\ : InMux
    port map (
            O => \N__38459\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__8233\ : CascadeMux
    port map (
            O => \N__38456\,
            I => \N__38453\
        );

    \I__8232\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38448\
        );

    \I__8231\ : InMux
    port map (
            O => \N__38452\,
            I => \N__38445\
        );

    \I__8230\ : InMux
    port map (
            O => \N__38451\,
            I => \N__38442\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__38448\,
            I => \N__38437\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__38445\,
            I => \N__38437\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__38442\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__8226\ : Odrv4
    port map (
            O => \N__38437\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__8225\ : InMux
    port map (
            O => \N__38432\,
            I => \bfn_16_25_0_\
        );

    \I__8224\ : CascadeMux
    port map (
            O => \N__38429\,
            I => \N__38425\
        );

    \I__8223\ : CascadeMux
    port map (
            O => \N__38428\,
            I => \N__38422\
        );

    \I__8222\ : InMux
    port map (
            O => \N__38425\,
            I => \N__38418\
        );

    \I__8221\ : InMux
    port map (
            O => \N__38422\,
            I => \N__38415\
        );

    \I__8220\ : InMux
    port map (
            O => \N__38421\,
            I => \N__38412\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__38418\,
            I => \N__38407\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__38415\,
            I => \N__38407\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__38412\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__38407\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__8215\ : InMux
    port map (
            O => \N__38402\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__8214\ : InMux
    port map (
            O => \N__38399\,
            I => \N__38392\
        );

    \I__8213\ : InMux
    port map (
            O => \N__38398\,
            I => \N__38392\
        );

    \I__8212\ : InMux
    port map (
            O => \N__38397\,
            I => \N__38389\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__38392\,
            I => \N__38386\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__38389\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__8209\ : Odrv4
    port map (
            O => \N__38386\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__8208\ : InMux
    port map (
            O => \N__38381\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__8207\ : CascadeMux
    port map (
            O => \N__38378\,
            I => \N__38375\
        );

    \I__8206\ : InMux
    port map (
            O => \N__38375\,
            I => \N__38370\
        );

    \I__8205\ : InMux
    port map (
            O => \N__38374\,
            I => \N__38367\
        );

    \I__8204\ : InMux
    port map (
            O => \N__38373\,
            I => \N__38364\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__38370\,
            I => \N__38359\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__38367\,
            I => \N__38359\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__38364\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__38359\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__8199\ : InMux
    port map (
            O => \N__38354\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__8198\ : CascadeMux
    port map (
            O => \N__38351\,
            I => \N__38348\
        );

    \I__8197\ : InMux
    port map (
            O => \N__38348\,
            I => \N__38343\
        );

    \I__8196\ : InMux
    port map (
            O => \N__38347\,
            I => \N__38340\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38346\,
            I => \N__38337\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__38343\,
            I => \N__38332\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__38340\,
            I => \N__38332\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__38337\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__8191\ : Odrv4
    port map (
            O => \N__38332\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__8190\ : InMux
    port map (
            O => \N__38327\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__8189\ : CascadeMux
    port map (
            O => \N__38324\,
            I => \N__38320\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38323\,
            I => \N__38316\
        );

    \I__8187\ : InMux
    port map (
            O => \N__38320\,
            I => \N__38313\
        );

    \I__8186\ : InMux
    port map (
            O => \N__38319\,
            I => \N__38310\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38316\,
            I => \N__38305\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__38313\,
            I => \N__38305\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__38310\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__8182\ : Odrv4
    port map (
            O => \N__38305\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__8181\ : InMux
    port map (
            O => \N__38300\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__38297\,
            I => \N__38294\
        );

    \I__8179\ : InMux
    port map (
            O => \N__38294\,
            I => \N__38289\
        );

    \I__8178\ : InMux
    port map (
            O => \N__38293\,
            I => \N__38286\
        );

    \I__8177\ : InMux
    port map (
            O => \N__38292\,
            I => \N__38283\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__38289\,
            I => \N__38278\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__38286\,
            I => \N__38278\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__38283\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__8173\ : Odrv4
    port map (
            O => \N__38278\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38273\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__38270\,
            I => \N__38266\
        );

    \I__8170\ : CascadeMux
    port map (
            O => \N__38269\,
            I => \N__38263\
        );

    \I__8169\ : InMux
    port map (
            O => \N__38266\,
            I => \N__38257\
        );

    \I__8168\ : InMux
    port map (
            O => \N__38263\,
            I => \N__38257\
        );

    \I__8167\ : InMux
    port map (
            O => \N__38262\,
            I => \N__38254\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__38257\,
            I => \N__38251\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__38254\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__8164\ : Odrv4
    port map (
            O => \N__38251\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38246\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38243\,
            I => \N__38236\
        );

    \I__8161\ : InMux
    port map (
            O => \N__38242\,
            I => \N__38236\
        );

    \I__8160\ : InMux
    port map (
            O => \N__38241\,
            I => \N__38233\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__38236\,
            I => \N__38230\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__38233\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__38230\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__8156\ : InMux
    port map (
            O => \N__38225\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__8155\ : CascadeMux
    port map (
            O => \N__38222\,
            I => \N__38219\
        );

    \I__8154\ : InMux
    port map (
            O => \N__38219\,
            I => \N__38214\
        );

    \I__8153\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38211\
        );

    \I__8152\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38208\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__38214\,
            I => \N__38203\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__38211\,
            I => \N__38203\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__38208\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__8148\ : Odrv4
    port map (
            O => \N__38203\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__8147\ : InMux
    port map (
            O => \N__38198\,
            I => \bfn_16_24_0_\
        );

    \I__8146\ : CascadeMux
    port map (
            O => \N__38195\,
            I => \N__38191\
        );

    \I__8145\ : CascadeMux
    port map (
            O => \N__38194\,
            I => \N__38188\
        );

    \I__8144\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38185\
        );

    \I__8143\ : InMux
    port map (
            O => \N__38188\,
            I => \N__38181\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__38185\,
            I => \N__38178\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38184\,
            I => \N__38175\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__38181\,
            I => \N__38170\
        );

    \I__8139\ : Span4Mux_h
    port map (
            O => \N__38178\,
            I => \N__38170\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38175\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__8137\ : Odrv4
    port map (
            O => \N__38170\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__8136\ : InMux
    port map (
            O => \N__38165\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__8135\ : InMux
    port map (
            O => \N__38162\,
            I => \N__38155\
        );

    \I__8134\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38155\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38152\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__38155\,
            I => \N__38149\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__38152\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__8130\ : Odrv4
    port map (
            O => \N__38149\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38144\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__8128\ : CascadeMux
    port map (
            O => \N__38141\,
            I => \N__38138\
        );

    \I__8127\ : InMux
    port map (
            O => \N__38138\,
            I => \N__38133\
        );

    \I__8126\ : InMux
    port map (
            O => \N__38137\,
            I => \N__38130\
        );

    \I__8125\ : InMux
    port map (
            O => \N__38136\,
            I => \N__38127\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38133\,
            I => \N__38122\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__38130\,
            I => \N__38122\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__38127\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__8121\ : Odrv4
    port map (
            O => \N__38122\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__8120\ : CascadeMux
    port map (
            O => \N__38117\,
            I => \N__38114\
        );

    \I__8119\ : InMux
    port map (
            O => \N__38114\,
            I => \N__38109\
        );

    \I__8118\ : InMux
    port map (
            O => \N__38113\,
            I => \N__38106\
        );

    \I__8117\ : InMux
    port map (
            O => \N__38112\,
            I => \N__38103\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__38109\,
            I => \N__38098\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__38106\,
            I => \N__38098\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__38103\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__8113\ : Odrv4
    port map (
            O => \N__38098\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__8112\ : InMux
    port map (
            O => \N__38093\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__8111\ : InMux
    port map (
            O => \N__38090\,
            I => \N__38083\
        );

    \I__8110\ : InMux
    port map (
            O => \N__38089\,
            I => \N__38083\
        );

    \I__8109\ : InMux
    port map (
            O => \N__38088\,
            I => \N__38080\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__38083\,
            I => \N__38077\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__38080\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__38077\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__8105\ : InMux
    port map (
            O => \N__38072\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__8104\ : CascadeMux
    port map (
            O => \N__38069\,
            I => \N__38066\
        );

    \I__8103\ : InMux
    port map (
            O => \N__38066\,
            I => \N__38061\
        );

    \I__8102\ : InMux
    port map (
            O => \N__38065\,
            I => \N__38058\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38064\,
            I => \N__38055\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__38061\,
            I => \N__38050\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__38058\,
            I => \N__38050\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__38055\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__8097\ : Odrv4
    port map (
            O => \N__38050\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__8096\ : InMux
    port map (
            O => \N__38045\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__8095\ : CascadeMux
    port map (
            O => \N__38042\,
            I => \N__38038\
        );

    \I__8094\ : CascadeMux
    port map (
            O => \N__38041\,
            I => \N__38035\
        );

    \I__8093\ : InMux
    port map (
            O => \N__38038\,
            I => \N__38029\
        );

    \I__8092\ : InMux
    port map (
            O => \N__38035\,
            I => \N__38029\
        );

    \I__8091\ : InMux
    port map (
            O => \N__38034\,
            I => \N__38026\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__38029\,
            I => \N__38023\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__38026\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__8088\ : Odrv4
    port map (
            O => \N__38023\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__8087\ : InMux
    port map (
            O => \N__38018\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__8086\ : InMux
    port map (
            O => \N__38015\,
            I => \N__38008\
        );

    \I__8085\ : InMux
    port map (
            O => \N__38014\,
            I => \N__38008\
        );

    \I__8084\ : InMux
    port map (
            O => \N__38013\,
            I => \N__38005\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__38008\,
            I => \N__38002\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__38005\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__8081\ : Odrv4
    port map (
            O => \N__38002\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__8080\ : InMux
    port map (
            O => \N__37997\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__8079\ : CascadeMux
    port map (
            O => \N__37994\,
            I => \N__37991\
        );

    \I__8078\ : InMux
    port map (
            O => \N__37991\,
            I => \N__37986\
        );

    \I__8077\ : InMux
    port map (
            O => \N__37990\,
            I => \N__37983\
        );

    \I__8076\ : InMux
    port map (
            O => \N__37989\,
            I => \N__37980\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__37986\,
            I => \N__37975\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__37983\,
            I => \N__37975\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__37980\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__8072\ : Odrv4
    port map (
            O => \N__37975\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__8071\ : InMux
    port map (
            O => \N__37970\,
            I => \bfn_16_23_0_\
        );

    \I__8070\ : CascadeMux
    port map (
            O => \N__37967\,
            I => \N__37963\
        );

    \I__8069\ : CascadeMux
    port map (
            O => \N__37966\,
            I => \N__37960\
        );

    \I__8068\ : InMux
    port map (
            O => \N__37963\,
            I => \N__37956\
        );

    \I__8067\ : InMux
    port map (
            O => \N__37960\,
            I => \N__37953\
        );

    \I__8066\ : InMux
    port map (
            O => \N__37959\,
            I => \N__37950\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__37956\,
            I => \N__37945\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__37953\,
            I => \N__37945\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__37950\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__8062\ : Odrv4
    port map (
            O => \N__37945\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__8061\ : InMux
    port map (
            O => \N__37940\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__8060\ : InMux
    port map (
            O => \N__37937\,
            I => \N__37930\
        );

    \I__8059\ : InMux
    port map (
            O => \N__37936\,
            I => \N__37930\
        );

    \I__8058\ : InMux
    port map (
            O => \N__37935\,
            I => \N__37927\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__37930\,
            I => \N__37924\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__37927\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__8055\ : Odrv4
    port map (
            O => \N__37924\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__8054\ : InMux
    port map (
            O => \N__37919\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__8053\ : CascadeMux
    port map (
            O => \N__37916\,
            I => \N__37908\
        );

    \I__8052\ : CascadeMux
    port map (
            O => \N__37915\,
            I => \N__37904\
        );

    \I__8051\ : CascadeMux
    port map (
            O => \N__37914\,
            I => \N__37900\
        );

    \I__8050\ : CascadeMux
    port map (
            O => \N__37913\,
            I => \N__37892\
        );

    \I__8049\ : CascadeMux
    port map (
            O => \N__37912\,
            I => \N__37888\
        );

    \I__8048\ : InMux
    port map (
            O => \N__37911\,
            I => \N__37864\
        );

    \I__8047\ : InMux
    port map (
            O => \N__37908\,
            I => \N__37864\
        );

    \I__8046\ : InMux
    port map (
            O => \N__37907\,
            I => \N__37864\
        );

    \I__8045\ : InMux
    port map (
            O => \N__37904\,
            I => \N__37864\
        );

    \I__8044\ : InMux
    port map (
            O => \N__37903\,
            I => \N__37864\
        );

    \I__8043\ : InMux
    port map (
            O => \N__37900\,
            I => \N__37864\
        );

    \I__8042\ : InMux
    port map (
            O => \N__37899\,
            I => \N__37864\
        );

    \I__8041\ : InMux
    port map (
            O => \N__37898\,
            I => \N__37859\
        );

    \I__8040\ : InMux
    port map (
            O => \N__37897\,
            I => \N__37859\
        );

    \I__8039\ : InMux
    port map (
            O => \N__37896\,
            I => \N__37846\
        );

    \I__8038\ : InMux
    port map (
            O => \N__37895\,
            I => \N__37846\
        );

    \I__8037\ : InMux
    port map (
            O => \N__37892\,
            I => \N__37846\
        );

    \I__8036\ : InMux
    port map (
            O => \N__37891\,
            I => \N__37846\
        );

    \I__8035\ : InMux
    port map (
            O => \N__37888\,
            I => \N__37846\
        );

    \I__8034\ : InMux
    port map (
            O => \N__37887\,
            I => \N__37846\
        );

    \I__8033\ : CascadeMux
    port map (
            O => \N__37886\,
            I => \N__37843\
        );

    \I__8032\ : CascadeMux
    port map (
            O => \N__37885\,
            I => \N__37839\
        );

    \I__8031\ : CascadeMux
    port map (
            O => \N__37884\,
            I => \N__37835\
        );

    \I__8030\ : CascadeMux
    port map (
            O => \N__37883\,
            I => \N__37831\
        );

    \I__8029\ : CascadeMux
    port map (
            O => \N__37882\,
            I => \N__37826\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__37881\,
            I => \N__37822\
        );

    \I__8027\ : CascadeMux
    port map (
            O => \N__37880\,
            I => \N__37818\
        );

    \I__8026\ : InMux
    port map (
            O => \N__37879\,
            I => \N__37814\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__37864\,
            I => \N__37796\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__37859\,
            I => \N__37796\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__37846\,
            I => \N__37796\
        );

    \I__8022\ : InMux
    port map (
            O => \N__37843\,
            I => \N__37779\
        );

    \I__8021\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37779\
        );

    \I__8020\ : InMux
    port map (
            O => \N__37839\,
            I => \N__37779\
        );

    \I__8019\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37779\
        );

    \I__8018\ : InMux
    port map (
            O => \N__37835\,
            I => \N__37779\
        );

    \I__8017\ : InMux
    port map (
            O => \N__37834\,
            I => \N__37779\
        );

    \I__8016\ : InMux
    port map (
            O => \N__37831\,
            I => \N__37779\
        );

    \I__8015\ : InMux
    port map (
            O => \N__37830\,
            I => \N__37779\
        );

    \I__8014\ : InMux
    port map (
            O => \N__37829\,
            I => \N__37764\
        );

    \I__8013\ : InMux
    port map (
            O => \N__37826\,
            I => \N__37764\
        );

    \I__8012\ : InMux
    port map (
            O => \N__37825\,
            I => \N__37764\
        );

    \I__8011\ : InMux
    port map (
            O => \N__37822\,
            I => \N__37764\
        );

    \I__8010\ : InMux
    port map (
            O => \N__37821\,
            I => \N__37764\
        );

    \I__8009\ : InMux
    port map (
            O => \N__37818\,
            I => \N__37764\
        );

    \I__8008\ : InMux
    port map (
            O => \N__37817\,
            I => \N__37764\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__37814\,
            I => \N__37759\
        );

    \I__8006\ : InMux
    port map (
            O => \N__37813\,
            I => \N__37756\
        );

    \I__8005\ : InMux
    port map (
            O => \N__37812\,
            I => \N__37753\
        );

    \I__8004\ : InMux
    port map (
            O => \N__37811\,
            I => \N__37750\
        );

    \I__8003\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37747\
        );

    \I__8002\ : InMux
    port map (
            O => \N__37809\,
            I => \N__37740\
        );

    \I__8001\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37740\
        );

    \I__8000\ : InMux
    port map (
            O => \N__37807\,
            I => \N__37740\
        );

    \I__7999\ : InMux
    port map (
            O => \N__37806\,
            I => \N__37731\
        );

    \I__7998\ : InMux
    port map (
            O => \N__37805\,
            I => \N__37731\
        );

    \I__7997\ : InMux
    port map (
            O => \N__37804\,
            I => \N__37731\
        );

    \I__7996\ : InMux
    port map (
            O => \N__37803\,
            I => \N__37731\
        );

    \I__7995\ : Span4Mux_v
    port map (
            O => \N__37796\,
            I => \N__37715\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__37779\,
            I => \N__37715\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__37764\,
            I => \N__37715\
        );

    \I__7992\ : InMux
    port map (
            O => \N__37763\,
            I => \N__37710\
        );

    \I__7991\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37710\
        );

    \I__7990\ : Span12Mux_s2_h
    port map (
            O => \N__37759\,
            I => \N__37707\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__37756\,
            I => \N__37700\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__37753\,
            I => \N__37700\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__37750\,
            I => \N__37700\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__37747\,
            I => \N__37693\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__37740\,
            I => \N__37693\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__37731\,
            I => \N__37693\
        );

    \I__7983\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37690\
        );

    \I__7982\ : InMux
    port map (
            O => \N__37729\,
            I => \N__37683\
        );

    \I__7981\ : InMux
    port map (
            O => \N__37728\,
            I => \N__37683\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37727\,
            I => \N__37683\
        );

    \I__7979\ : InMux
    port map (
            O => \N__37726\,
            I => \N__37674\
        );

    \I__7978\ : InMux
    port map (
            O => \N__37725\,
            I => \N__37674\
        );

    \I__7977\ : InMux
    port map (
            O => \N__37724\,
            I => \N__37674\
        );

    \I__7976\ : InMux
    port map (
            O => \N__37723\,
            I => \N__37674\
        );

    \I__7975\ : CascadeMux
    port map (
            O => \N__37722\,
            I => \N__37670\
        );

    \I__7974\ : Span4Mux_v
    port map (
            O => \N__37715\,
            I => \N__37664\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__37710\,
            I => \N__37664\
        );

    \I__7972\ : Span12Mux_v
    port map (
            O => \N__37707\,
            I => \N__37661\
        );

    \I__7971\ : Span12Mux_s8_v
    port map (
            O => \N__37700\,
            I => \N__37650\
        );

    \I__7970\ : Span12Mux_s9_v
    port map (
            O => \N__37693\,
            I => \N__37650\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__37690\,
            I => \N__37650\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__37683\,
            I => \N__37650\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__37674\,
            I => \N__37650\
        );

    \I__7966\ : InMux
    port map (
            O => \N__37673\,
            I => \N__37643\
        );

    \I__7965\ : InMux
    port map (
            O => \N__37670\,
            I => \N__37643\
        );

    \I__7964\ : InMux
    port map (
            O => \N__37669\,
            I => \N__37643\
        );

    \I__7963\ : Span4Mux_v
    port map (
            O => \N__37664\,
            I => \N__37640\
        );

    \I__7962\ : Span12Mux_h
    port map (
            O => \N__37661\,
            I => \N__37637\
        );

    \I__7961\ : Span12Mux_v
    port map (
            O => \N__37650\,
            I => \N__37632\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__37643\,
            I => \N__37632\
        );

    \I__7959\ : Span4Mux_h
    port map (
            O => \N__37640\,
            I => \N__37629\
        );

    \I__7958\ : Odrv12
    port map (
            O => \N__37637\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7957\ : Odrv12
    port map (
            O => \N__37632\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7956\ : Odrv4
    port map (
            O => \N__37629\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7955\ : CascadeMux
    port map (
            O => \N__37622\,
            I => \N__37619\
        );

    \I__7954\ : InMux
    port map (
            O => \N__37619\,
            I => \N__37616\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__37616\,
            I => \N__37613\
        );

    \I__7952\ : Span4Mux_h
    port map (
            O => \N__37613\,
            I => \N__37610\
        );

    \I__7951\ : Odrv4
    port map (
            O => \N__37610\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__7950\ : InMux
    port map (
            O => \N__37607\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__7949\ : InMux
    port map (
            O => \N__37604\,
            I => \N__37601\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__37601\,
            I => \N__37598\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__37598\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__7946\ : CascadeMux
    port map (
            O => \N__37595\,
            I => \N__37592\
        );

    \I__7945\ : InMux
    port map (
            O => \N__37592\,
            I => \N__37589\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__37589\,
            I => \N__37586\
        );

    \I__7943\ : Odrv4
    port map (
            O => \N__37586\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__7942\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37580\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__37580\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__7940\ : InMux
    port map (
            O => \N__37577\,
            I => \N__37574\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__37574\,
            I => \N__37571\
        );

    \I__7938\ : Span4Mux_h
    port map (
            O => \N__37571\,
            I => \N__37568\
        );

    \I__7937\ : Odrv4
    port map (
            O => \N__37568\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__7936\ : InMux
    port map (
            O => \N__37565\,
            I => \N__37562\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__37562\,
            I => \N__37559\
        );

    \I__7934\ : Span4Mux_v
    port map (
            O => \N__37559\,
            I => \N__37555\
        );

    \I__7933\ : InMux
    port map (
            O => \N__37558\,
            I => \N__37551\
        );

    \I__7932\ : Span4Mux_h
    port map (
            O => \N__37555\,
            I => \N__37548\
        );

    \I__7931\ : InMux
    port map (
            O => \N__37554\,
            I => \N__37545\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__37551\,
            I => \N__37542\
        );

    \I__7929\ : Odrv4
    port map (
            O => \N__37548\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__37545\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__7927\ : Odrv4
    port map (
            O => \N__37542\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__7926\ : InMux
    port map (
            O => \N__37535\,
            I => \bfn_16_22_0_\
        );

    \I__7925\ : InMux
    port map (
            O => \N__37532\,
            I => \N__37529\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__37529\,
            I => \N__37525\
        );

    \I__7923\ : CascadeMux
    port map (
            O => \N__37528\,
            I => \N__37522\
        );

    \I__7922\ : Span4Mux_v
    port map (
            O => \N__37525\,
            I => \N__37519\
        );

    \I__7921\ : InMux
    port map (
            O => \N__37522\,
            I => \N__37515\
        );

    \I__7920\ : Span4Mux_h
    port map (
            O => \N__37519\,
            I => \N__37512\
        );

    \I__7919\ : InMux
    port map (
            O => \N__37518\,
            I => \N__37509\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__37515\,
            I => \N__37506\
        );

    \I__7917\ : Odrv4
    port map (
            O => \N__37512\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__37509\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__7915\ : Odrv4
    port map (
            O => \N__37506\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__7914\ : InMux
    port map (
            O => \N__37499\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__7913\ : CascadeMux
    port map (
            O => \N__37496\,
            I => \N__37492\
        );

    \I__7912\ : CascadeMux
    port map (
            O => \N__37495\,
            I => \N__37489\
        );

    \I__7911\ : InMux
    port map (
            O => \N__37492\,
            I => \N__37484\
        );

    \I__7910\ : InMux
    port map (
            O => \N__37489\,
            I => \N__37484\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__37484\,
            I => \N__37480\
        );

    \I__7908\ : InMux
    port map (
            O => \N__37483\,
            I => \N__37477\
        );

    \I__7907\ : Span12Mux_h
    port map (
            O => \N__37480\,
            I => \N__37474\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__37477\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__7905\ : Odrv12
    port map (
            O => \N__37474\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__7904\ : InMux
    port map (
            O => \N__37469\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__7903\ : CascadeMux
    port map (
            O => \N__37466\,
            I => \N__37463\
        );

    \I__7902\ : InMux
    port map (
            O => \N__37463\,
            I => \N__37460\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__37460\,
            I => \N__37457\
        );

    \I__7900\ : Span4Mux_v
    port map (
            O => \N__37457\,
            I => \N__37454\
        );

    \I__7899\ : Span4Mux_h
    port map (
            O => \N__37454\,
            I => \N__37451\
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__37451\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__7897\ : InMux
    port map (
            O => \N__37448\,
            I => \N__37445\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__37445\,
            I => \N__37442\
        );

    \I__7895\ : Span4Mux_h
    port map (
            O => \N__37442\,
            I => \N__37439\
        );

    \I__7894\ : Span4Mux_v
    port map (
            O => \N__37439\,
            I => \N__37436\
        );

    \I__7893\ : Odrv4
    port map (
            O => \N__37436\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__7892\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37430\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__37430\,
            I => \N__37427\
        );

    \I__7890\ : Span4Mux_h
    port map (
            O => \N__37427\,
            I => \N__37424\
        );

    \I__7889\ : Odrv4
    port map (
            O => \N__37424\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__7888\ : CascadeMux
    port map (
            O => \N__37421\,
            I => \N__37418\
        );

    \I__7887\ : InMux
    port map (
            O => \N__37418\,
            I => \N__37415\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__37415\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__7885\ : InMux
    port map (
            O => \N__37412\,
            I => \N__37409\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__37409\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__7883\ : CascadeMux
    port map (
            O => \N__37406\,
            I => \N__37403\
        );

    \I__7882\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37400\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__37400\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__7880\ : CascadeMux
    port map (
            O => \N__37397\,
            I => \N__37394\
        );

    \I__7879\ : InMux
    port map (
            O => \N__37394\,
            I => \N__37391\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__37391\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__7877\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37385\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__37385\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__7875\ : CascadeMux
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__7874\ : InMux
    port map (
            O => \N__37379\,
            I => \N__37376\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__37376\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__7872\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37370\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__37370\,
            I => \N__37367\
        );

    \I__7870\ : Span4Mux_h
    port map (
            O => \N__37367\,
            I => \N__37364\
        );

    \I__7869\ : Odrv4
    port map (
            O => \N__37364\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__7868\ : CascadeMux
    port map (
            O => \N__37361\,
            I => \N__37358\
        );

    \I__7867\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37355\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__37355\,
            I => \N__37352\
        );

    \I__7865\ : Span12Mux_v
    port map (
            O => \N__37352\,
            I => \N__37349\
        );

    \I__7864\ : Odrv12
    port map (
            O => \N__37349\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__7863\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37343\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__37343\,
            I => \N__37340\
        );

    \I__7861\ : Span4Mux_v
    port map (
            O => \N__37340\,
            I => \N__37337\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__37337\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__7859\ : CascadeMux
    port map (
            O => \N__37334\,
            I => \N__37331\
        );

    \I__7858\ : InMux
    port map (
            O => \N__37331\,
            I => \N__37328\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__37328\,
            I => \N__37325\
        );

    \I__7856\ : Span4Mux_h
    port map (
            O => \N__37325\,
            I => \N__37322\
        );

    \I__7855\ : Odrv4
    port map (
            O => \N__37322\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__7854\ : InMux
    port map (
            O => \N__37319\,
            I => \N__37316\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__37316\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__7852\ : CascadeMux
    port map (
            O => \N__37313\,
            I => \N__37310\
        );

    \I__7851\ : InMux
    port map (
            O => \N__37310\,
            I => \N__37307\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__37307\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37304\,
            I => \N__37301\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__37301\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37298\,
            I => \N__37295\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__37295\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__7845\ : CascadeMux
    port map (
            O => \N__37292\,
            I => \N__37289\
        );

    \I__7844\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37286\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__37286\,
            I => \current_shift_inst.control_input_1_axb_1\
        );

    \I__7842\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37280\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__37280\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37274\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__37274\,
            I => \current_shift_inst.control_input_1_axb_7\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37271\,
            I => \N__37268\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__37268\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__7836\ : InMux
    port map (
            O => \N__37265\,
            I => \N__37262\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__37262\,
            I => \current_shift_inst.control_input_1_axb_10\
        );

    \I__7834\ : InMux
    port map (
            O => \N__37259\,
            I => \N__37256\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__37256\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__7832\ : InMux
    port map (
            O => \N__37253\,
            I => \N__37250\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__37250\,
            I => \current_shift_inst.control_input_1_axb_2\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37247\,
            I => \N__37244\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__37244\,
            I => \N__37241\
        );

    \I__7828\ : Span4Mux_h
    port map (
            O => \N__37241\,
            I => \N__37237\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37240\,
            I => \N__37234\
        );

    \I__7826\ : Span4Mux_v
    port map (
            O => \N__37237\,
            I => \N__37231\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__37234\,
            I => \N__37228\
        );

    \I__7824\ : Odrv4
    port map (
            O => \N__37231\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__7823\ : Odrv12
    port map (
            O => \N__37228\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__7822\ : CascadeMux
    port map (
            O => \N__37223\,
            I => \N__37220\
        );

    \I__7821\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37217\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__37217\,
            I => \N__37212\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37216\,
            I => \N__37207\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37215\,
            I => \N__37207\
        );

    \I__7817\ : Odrv12
    port map (
            O => \N__37212\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__37207\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__7815\ : CascadeMux
    port map (
            O => \N__37202\,
            I => \N__37199\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37199\,
            I => \N__37196\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__37196\,
            I => \N__37193\
        );

    \I__7812\ : Odrv12
    port map (
            O => \N__37193\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__7811\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37187\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__37187\,
            I => \N__37184\
        );

    \I__7809\ : Span4Mux_h
    port map (
            O => \N__37184\,
            I => \N__37181\
        );

    \I__7808\ : Odrv4
    port map (
            O => \N__37181\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__7807\ : CascadeMux
    port map (
            O => \N__37178\,
            I => \N__37175\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37175\,
            I => \N__37172\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__37172\,
            I => \N__37169\
        );

    \I__7804\ : Odrv4
    port map (
            O => \N__37169\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37166\,
            I => \N__37163\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__37163\,
            I => \N__37160\
        );

    \I__7801\ : Odrv12
    port map (
            O => \N__37160\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__7800\ : InMux
    port map (
            O => \N__37157\,
            I => \current_shift_inst.control_input_1_cry_2\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37154\,
            I => \N__37151\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__37151\,
            I => \current_shift_inst.control_input_1_axb_4\
        );

    \I__7797\ : InMux
    port map (
            O => \N__37148\,
            I => \N__37145\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__37145\,
            I => \N__37142\
        );

    \I__7795\ : Span12Mux_v
    port map (
            O => \N__37142\,
            I => \N__37139\
        );

    \I__7794\ : Odrv12
    port map (
            O => \N__37139\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__7793\ : InMux
    port map (
            O => \N__37136\,
            I => \current_shift_inst.control_input_1_cry_3\
        );

    \I__7792\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37130\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__37130\,
            I => \current_shift_inst.control_input_1_axb_5\
        );

    \I__7790\ : InMux
    port map (
            O => \N__37127\,
            I => \N__37124\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__37124\,
            I => \N__37121\
        );

    \I__7788\ : Span4Mux_v
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__7787\ : Span4Mux_h
    port map (
            O => \N__37118\,
            I => \N__37115\
        );

    \I__7786\ : Odrv4
    port map (
            O => \N__37115\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__7785\ : InMux
    port map (
            O => \N__37112\,
            I => \current_shift_inst.control_input_1_cry_4\
        );

    \I__7784\ : InMux
    port map (
            O => \N__37109\,
            I => \N__37106\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__37106\,
            I => \N__37103\
        );

    \I__7782\ : Odrv12
    port map (
            O => \N__37103\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__7781\ : InMux
    port map (
            O => \N__37100\,
            I => \current_shift_inst.control_input_1_cry_5\
        );

    \I__7780\ : InMux
    port map (
            O => \N__37097\,
            I => \N__37094\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__37094\,
            I => \N__37091\
        );

    \I__7778\ : Span4Mux_h
    port map (
            O => \N__37091\,
            I => \N__37088\
        );

    \I__7777\ : Span4Mux_h
    port map (
            O => \N__37088\,
            I => \N__37085\
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__37085\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__7775\ : InMux
    port map (
            O => \N__37082\,
            I => \current_shift_inst.control_input_1_cry_6\
        );

    \I__7774\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37076\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__37076\,
            I => \N__37073\
        );

    \I__7772\ : Span4Mux_h
    port map (
            O => \N__37073\,
            I => \N__37070\
        );

    \I__7771\ : Odrv4
    port map (
            O => \N__37070\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__7770\ : InMux
    port map (
            O => \N__37067\,
            I => \bfn_16_16_0_\
        );

    \I__7769\ : InMux
    port map (
            O => \N__37064\,
            I => \current_shift_inst.control_input_1_cry_8\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37061\,
            I => \N__37058\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__37058\,
            I => \N__37055\
        );

    \I__7766\ : Span4Mux_v
    port map (
            O => \N__37055\,
            I => \N__37052\
        );

    \I__7765\ : Odrv4
    port map (
            O => \N__37052\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__7764\ : InMux
    port map (
            O => \N__37049\,
            I => \current_shift_inst.control_input_1_cry_9\
        );

    \I__7763\ : InMux
    port map (
            O => \N__37046\,
            I => \N__37043\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__37043\,
            I => \current_shift_inst.control_input_1_axb_11\
        );

    \I__7761\ : InMux
    port map (
            O => \N__37040\,
            I => \current_shift_inst.control_input_1_cry_10\
        );

    \I__7760\ : InMux
    port map (
            O => \N__37037\,
            I => \N__37034\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__37034\,
            I => \N__37030\
        );

    \I__7758\ : InMux
    port map (
            O => \N__37033\,
            I => \N__37027\
        );

    \I__7757\ : Span12Mux_s9_h
    port map (
            O => \N__37030\,
            I => \N__37024\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__37027\,
            I => \N__37021\
        );

    \I__7755\ : Odrv12
    port map (
            O => \N__37024\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__7754\ : Odrv4
    port map (
            O => \N__37021\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__7753\ : InMux
    port map (
            O => \N__37016\,
            I => \N__37013\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__7751\ : Odrv4
    port map (
            O => \N__37010\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__7750\ : InMux
    port map (
            O => \N__37007\,
            I => \N__37004\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__37004\,
            I => \N__37001\
        );

    \I__7748\ : Odrv4
    port map (
            O => \N__37001\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__7747\ : InMux
    port map (
            O => \N__36998\,
            I => \N__36995\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__36995\,
            I => \N__36992\
        );

    \I__7745\ : Span12Mux_v
    port map (
            O => \N__36992\,
            I => \N__36989\
        );

    \I__7744\ : Odrv12
    port map (
            O => \N__36989\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__7743\ : CascadeMux
    port map (
            O => \N__36986\,
            I => \N__36982\
        );

    \I__7742\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36978\
        );

    \I__7741\ : InMux
    port map (
            O => \N__36982\,
            I => \N__36975\
        );

    \I__7740\ : InMux
    port map (
            O => \N__36981\,
            I => \N__36972\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__36978\,
            I => \N__36969\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__36975\,
            I => \N__36966\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__36972\,
            I => \N__36963\
        );

    \I__7736\ : Span4Mux_h
    port map (
            O => \N__36969\,
            I => \N__36960\
        );

    \I__7735\ : Span4Mux_v
    port map (
            O => \N__36966\,
            I => \N__36955\
        );

    \I__7734\ : Span4Mux_h
    port map (
            O => \N__36963\,
            I => \N__36955\
        );

    \I__7733\ : Odrv4
    port map (
            O => \N__36960\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__7732\ : Odrv4
    port map (
            O => \N__36955\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__7731\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36947\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__36947\,
            I => \N__36944\
        );

    \I__7729\ : Odrv4
    port map (
            O => \N__36944\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__7728\ : InMux
    port map (
            O => \N__36941\,
            I => \N__36938\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__36938\,
            I => \current_shift_inst.control_input_1_axb_0\
        );

    \I__7726\ : InMux
    port map (
            O => \N__36935\,
            I => \N__36931\
        );

    \I__7725\ : CascadeMux
    port map (
            O => \N__36934\,
            I => \N__36928\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__36931\,
            I => \N__36925\
        );

    \I__7723\ : InMux
    port map (
            O => \N__36928\,
            I => \N__36922\
        );

    \I__7722\ : Odrv4
    port map (
            O => \N__36925\,
            I => \current_shift_inst.N_1572_i\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__36922\,
            I => \current_shift_inst.N_1572_i\
        );

    \I__7720\ : InMux
    port map (
            O => \N__36917\,
            I => \N__36913\
        );

    \I__7719\ : InMux
    port map (
            O => \N__36916\,
            I => \N__36910\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__36913\,
            I => \N__36905\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__36910\,
            I => \N__36905\
        );

    \I__7716\ : Span12Mux_h
    port map (
            O => \N__36905\,
            I => \N__36902\
        );

    \I__7715\ : Odrv12
    port map (
            O => \N__36902\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__7714\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36896\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__36896\,
            I => \N__36893\
        );

    \I__7712\ : Span4Mux_h
    port map (
            O => \N__36893\,
            I => \N__36890\
        );

    \I__7711\ : Span4Mux_h
    port map (
            O => \N__36890\,
            I => \N__36887\
        );

    \I__7710\ : Span4Mux_h
    port map (
            O => \N__36887\,
            I => \N__36884\
        );

    \I__7709\ : Odrv4
    port map (
            O => \N__36884\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__7708\ : InMux
    port map (
            O => \N__36881\,
            I => \current_shift_inst.control_input_1_cry_0\
        );

    \I__7707\ : InMux
    port map (
            O => \N__36878\,
            I => \N__36875\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__36875\,
            I => \N__36872\
        );

    \I__7705\ : Span4Mux_v
    port map (
            O => \N__36872\,
            I => \N__36869\
        );

    \I__7704\ : Span4Mux_h
    port map (
            O => \N__36869\,
            I => \N__36866\
        );

    \I__7703\ : Odrv4
    port map (
            O => \N__36866\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__7702\ : InMux
    port map (
            O => \N__36863\,
            I => \current_shift_inst.control_input_1_cry_1\
        );

    \I__7701\ : InMux
    port map (
            O => \N__36860\,
            I => \N__36857\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__36857\,
            I => \current_shift_inst.control_input_1_axb_3\
        );

    \I__7699\ : InMux
    port map (
            O => \N__36854\,
            I => \N__36850\
        );

    \I__7698\ : InMux
    port map (
            O => \N__36853\,
            I => \N__36847\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__36850\,
            I => \N__36844\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__36847\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__7695\ : Odrv4
    port map (
            O => \N__36844\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__7694\ : CascadeMux
    port map (
            O => \N__36839\,
            I => \N__36836\
        );

    \I__7693\ : InMux
    port map (
            O => \N__36836\,
            I => \N__36831\
        );

    \I__7692\ : InMux
    port map (
            O => \N__36835\,
            I => \N__36828\
        );

    \I__7691\ : InMux
    port map (
            O => \N__36834\,
            I => \N__36825\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__36831\,
            I => \N__36820\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__36828\,
            I => \N__36820\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__36825\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__7687\ : Odrv4
    port map (
            O => \N__36820\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__7686\ : InMux
    port map (
            O => \N__36815\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__7685\ : InMux
    port map (
            O => \N__36812\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__7684\ : IoInMux
    port map (
            O => \N__36809\,
            I => \N__36806\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__36806\,
            I => \N__36803\
        );

    \I__7682\ : Span12Mux_s8_v
    port map (
            O => \N__36803\,
            I => \N__36799\
        );

    \I__7681\ : InMux
    port map (
            O => \N__36802\,
            I => \N__36796\
        );

    \I__7680\ : Odrv12
    port map (
            O => \N__36799\,
            I => \T45_c\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__36796\,
            I => \T45_c\
        );

    \I__7678\ : CascadeMux
    port map (
            O => \N__36791\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__7677\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36785\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__36785\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__7675\ : InMux
    port map (
            O => \N__36782\,
            I => \N__36779\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__36779\,
            I => \N__36776\
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__36776\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__36773\,
            I => \N__36769\
        );

    \I__7671\ : InMux
    port map (
            O => \N__36772\,
            I => \N__36765\
        );

    \I__7670\ : InMux
    port map (
            O => \N__36769\,
            I => \N__36762\
        );

    \I__7669\ : InMux
    port map (
            O => \N__36768\,
            I => \N__36759\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__36765\,
            I => \N__36756\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__36762\,
            I => \N__36751\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__36759\,
            I => \N__36751\
        );

    \I__7665\ : Span4Mux_v
    port map (
            O => \N__36756\,
            I => \N__36747\
        );

    \I__7664\ : Span4Mux_h
    port map (
            O => \N__36751\,
            I => \N__36744\
        );

    \I__7663\ : InMux
    port map (
            O => \N__36750\,
            I => \N__36741\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__36747\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__7661\ : Odrv4
    port map (
            O => \N__36744\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__36741\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__7659\ : InMux
    port map (
            O => \N__36734\,
            I => \N__36731\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__36731\,
            I => \N__36728\
        );

    \I__7657\ : Span4Mux_v
    port map (
            O => \N__36728\,
            I => \N__36723\
        );

    \I__7656\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36718\
        );

    \I__7655\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36718\
        );

    \I__7654\ : Odrv4
    port map (
            O => \N__36723\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__36718\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__7652\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36706\
        );

    \I__7651\ : InMux
    port map (
            O => \N__36712\,
            I => \N__36706\
        );

    \I__7650\ : InMux
    port map (
            O => \N__36711\,
            I => \N__36703\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__36706\,
            I => \N__36700\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__36703\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__7647\ : Odrv4
    port map (
            O => \N__36700\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__7646\ : InMux
    port map (
            O => \N__36695\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__7645\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36685\
        );

    \I__7644\ : InMux
    port map (
            O => \N__36691\,
            I => \N__36685\
        );

    \I__7643\ : InMux
    port map (
            O => \N__36690\,
            I => \N__36682\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__36685\,
            I => \N__36679\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__36682\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__7640\ : Odrv4
    port map (
            O => \N__36679\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__7639\ : InMux
    port map (
            O => \N__36674\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__7638\ : CascadeMux
    port map (
            O => \N__36671\,
            I => \N__36667\
        );

    \I__7637\ : InMux
    port map (
            O => \N__36670\,
            I => \N__36663\
        );

    \I__7636\ : InMux
    port map (
            O => \N__36667\,
            I => \N__36660\
        );

    \I__7635\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36657\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__36663\,
            I => \N__36652\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__36660\,
            I => \N__36652\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__36657\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__7631\ : Odrv4
    port map (
            O => \N__36652\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__7630\ : InMux
    port map (
            O => \N__36647\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__7629\ : CascadeMux
    port map (
            O => \N__36644\,
            I => \N__36640\
        );

    \I__7628\ : InMux
    port map (
            O => \N__36643\,
            I => \N__36636\
        );

    \I__7627\ : InMux
    port map (
            O => \N__36640\,
            I => \N__36633\
        );

    \I__7626\ : InMux
    port map (
            O => \N__36639\,
            I => \N__36630\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__36636\,
            I => \N__36625\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__36633\,
            I => \N__36625\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__36630\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__7622\ : Odrv4
    port map (
            O => \N__36625\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__7621\ : InMux
    port map (
            O => \N__36620\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__7620\ : CascadeMux
    port map (
            O => \N__36617\,
            I => \N__36613\
        );

    \I__7619\ : CascadeMux
    port map (
            O => \N__36616\,
            I => \N__36610\
        );

    \I__7618\ : InMux
    port map (
            O => \N__36613\,
            I => \N__36604\
        );

    \I__7617\ : InMux
    port map (
            O => \N__36610\,
            I => \N__36604\
        );

    \I__7616\ : InMux
    port map (
            O => \N__36609\,
            I => \N__36601\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__36604\,
            I => \N__36598\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__36601\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__7613\ : Odrv4
    port map (
            O => \N__36598\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__7612\ : InMux
    port map (
            O => \N__36593\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__7611\ : CascadeMux
    port map (
            O => \N__36590\,
            I => \N__36586\
        );

    \I__7610\ : CascadeMux
    port map (
            O => \N__36589\,
            I => \N__36583\
        );

    \I__7609\ : InMux
    port map (
            O => \N__36586\,
            I => \N__36577\
        );

    \I__7608\ : InMux
    port map (
            O => \N__36583\,
            I => \N__36577\
        );

    \I__7607\ : InMux
    port map (
            O => \N__36582\,
            I => \N__36574\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__36577\,
            I => \N__36571\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__36574\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__7604\ : Odrv4
    port map (
            O => \N__36571\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__7603\ : InMux
    port map (
            O => \N__36566\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__7602\ : CascadeMux
    port map (
            O => \N__36563\,
            I => \N__36560\
        );

    \I__7601\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36557\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__36557\,
            I => \N__36552\
        );

    \I__7599\ : InMux
    port map (
            O => \N__36556\,
            I => \N__36549\
        );

    \I__7598\ : InMux
    port map (
            O => \N__36555\,
            I => \N__36546\
        );

    \I__7597\ : Span4Mux_v
    port map (
            O => \N__36552\,
            I => \N__36543\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__36549\,
            I => \N__36540\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__36546\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7594\ : Odrv4
    port map (
            O => \N__36543\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7593\ : Odrv4
    port map (
            O => \N__36540\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7592\ : InMux
    port map (
            O => \N__36533\,
            I => \bfn_16_11_0_\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__36530\,
            I => \N__36527\
        );

    \I__7590\ : InMux
    port map (
            O => \N__36527\,
            I => \N__36524\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__36524\,
            I => \N__36519\
        );

    \I__7588\ : InMux
    port map (
            O => \N__36523\,
            I => \N__36516\
        );

    \I__7587\ : InMux
    port map (
            O => \N__36522\,
            I => \N__36513\
        );

    \I__7586\ : Span4Mux_v
    port map (
            O => \N__36519\,
            I => \N__36508\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__36516\,
            I => \N__36508\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__36513\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__7583\ : Odrv4
    port map (
            O => \N__36508\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__7582\ : InMux
    port map (
            O => \N__36503\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__7581\ : InMux
    port map (
            O => \N__36500\,
            I => \N__36493\
        );

    \I__7580\ : InMux
    port map (
            O => \N__36499\,
            I => \N__36493\
        );

    \I__7579\ : InMux
    port map (
            O => \N__36498\,
            I => \N__36490\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__36493\,
            I => \N__36487\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__36490\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__7576\ : Odrv4
    port map (
            O => \N__36487\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__7575\ : CascadeMux
    port map (
            O => \N__36482\,
            I => \N__36479\
        );

    \I__7574\ : InMux
    port map (
            O => \N__36479\,
            I => \N__36476\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__36476\,
            I => \N__36472\
        );

    \I__7572\ : InMux
    port map (
            O => \N__36475\,
            I => \N__36469\
        );

    \I__7571\ : Span4Mux_h
    port map (
            O => \N__36472\,
            I => \N__36466\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__36469\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__7569\ : Odrv4
    port map (
            O => \N__36466\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__7568\ : InMux
    port map (
            O => \N__36461\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__7567\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36451\
        );

    \I__7566\ : InMux
    port map (
            O => \N__36457\,
            I => \N__36451\
        );

    \I__7565\ : InMux
    port map (
            O => \N__36456\,
            I => \N__36448\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__36451\,
            I => \N__36445\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__36448\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__7562\ : Odrv4
    port map (
            O => \N__36445\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__7561\ : InMux
    port map (
            O => \N__36440\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__7560\ : CascadeMux
    port map (
            O => \N__36437\,
            I => \N__36434\
        );

    \I__7559\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36429\
        );

    \I__7558\ : InMux
    port map (
            O => \N__36433\,
            I => \N__36426\
        );

    \I__7557\ : InMux
    port map (
            O => \N__36432\,
            I => \N__36423\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__36429\,
            I => \N__36418\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__36426\,
            I => \N__36418\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__36423\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__7553\ : Odrv4
    port map (
            O => \N__36418\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__7552\ : InMux
    port map (
            O => \N__36413\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__7551\ : CascadeMux
    port map (
            O => \N__36410\,
            I => \N__36406\
        );

    \I__7550\ : InMux
    port map (
            O => \N__36409\,
            I => \N__36402\
        );

    \I__7549\ : InMux
    port map (
            O => \N__36406\,
            I => \N__36399\
        );

    \I__7548\ : InMux
    port map (
            O => \N__36405\,
            I => \N__36396\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__36402\,
            I => \N__36391\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__36399\,
            I => \N__36391\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__36396\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__36391\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__7543\ : InMux
    port map (
            O => \N__36386\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__7542\ : InMux
    port map (
            O => \N__36383\,
            I => \N__36376\
        );

    \I__7541\ : InMux
    port map (
            O => \N__36382\,
            I => \N__36376\
        );

    \I__7540\ : InMux
    port map (
            O => \N__36381\,
            I => \N__36373\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__36376\,
            I => \N__36370\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__36373\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__7537\ : Odrv4
    port map (
            O => \N__36370\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__7536\ : InMux
    port map (
            O => \N__36365\,
            I => \N__36360\
        );

    \I__7535\ : InMux
    port map (
            O => \N__36364\,
            I => \N__36355\
        );

    \I__7534\ : InMux
    port map (
            O => \N__36363\,
            I => \N__36355\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__36360\,
            I => \N__36352\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__36355\,
            I => \N__36349\
        );

    \I__7531\ : Odrv4
    port map (
            O => \N__36352\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__7530\ : Odrv4
    port map (
            O => \N__36349\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__7529\ : InMux
    port map (
            O => \N__36344\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__7528\ : CascadeMux
    port map (
            O => \N__36341\,
            I => \N__36337\
        );

    \I__7527\ : CascadeMux
    port map (
            O => \N__36340\,
            I => \N__36334\
        );

    \I__7526\ : InMux
    port map (
            O => \N__36337\,
            I => \N__36328\
        );

    \I__7525\ : InMux
    port map (
            O => \N__36334\,
            I => \N__36328\
        );

    \I__7524\ : InMux
    port map (
            O => \N__36333\,
            I => \N__36325\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__36328\,
            I => \N__36322\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__36325\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__7521\ : Odrv4
    port map (
            O => \N__36322\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__7520\ : CascadeMux
    port map (
            O => \N__36317\,
            I => \N__36313\
        );

    \I__7519\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36310\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36313\,
            I => \N__36306\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__36310\,
            I => \N__36303\
        );

    \I__7516\ : InMux
    port map (
            O => \N__36309\,
            I => \N__36300\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__36306\,
            I => \N__36297\
        );

    \I__7514\ : Span4Mux_h
    port map (
            O => \N__36303\,
            I => \N__36292\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__36300\,
            I => \N__36292\
        );

    \I__7512\ : Odrv12
    port map (
            O => \N__36297\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__7511\ : Odrv4
    port map (
            O => \N__36292\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__7510\ : InMux
    port map (
            O => \N__36287\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__7509\ : CascadeMux
    port map (
            O => \N__36284\,
            I => \N__36280\
        );

    \I__7508\ : CascadeMux
    port map (
            O => \N__36283\,
            I => \N__36277\
        );

    \I__7507\ : InMux
    port map (
            O => \N__36280\,
            I => \N__36272\
        );

    \I__7506\ : InMux
    port map (
            O => \N__36277\,
            I => \N__36272\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__36272\,
            I => \N__36268\
        );

    \I__7504\ : InMux
    port map (
            O => \N__36271\,
            I => \N__36265\
        );

    \I__7503\ : Span4Mux_v
    port map (
            O => \N__36268\,
            I => \N__36262\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__36265\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__7501\ : Odrv4
    port map (
            O => \N__36262\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__7500\ : InMux
    port map (
            O => \N__36257\,
            I => \N__36254\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__36254\,
            I => \N__36249\
        );

    \I__7498\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36244\
        );

    \I__7497\ : InMux
    port map (
            O => \N__36252\,
            I => \N__36244\
        );

    \I__7496\ : Span4Mux_h
    port map (
            O => \N__36249\,
            I => \N__36239\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__36244\,
            I => \N__36239\
        );

    \I__7494\ : Odrv4
    port map (
            O => \N__36239\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__7493\ : InMux
    port map (
            O => \N__36236\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__7492\ : CascadeMux
    port map (
            O => \N__36233\,
            I => \N__36230\
        );

    \I__7491\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36227\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__36227\,
            I => \N__36222\
        );

    \I__7489\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36219\
        );

    \I__7488\ : InMux
    port map (
            O => \N__36225\,
            I => \N__36216\
        );

    \I__7487\ : Span4Mux_v
    port map (
            O => \N__36222\,
            I => \N__36211\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__36219\,
            I => \N__36211\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__36216\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__7484\ : Odrv4
    port map (
            O => \N__36211\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__7483\ : CascadeMux
    port map (
            O => \N__36206\,
            I => \N__36203\
        );

    \I__7482\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36200\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__36200\,
            I => \N__36195\
        );

    \I__7480\ : InMux
    port map (
            O => \N__36199\,
            I => \N__36190\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36190\
        );

    \I__7478\ : Span4Mux_v
    port map (
            O => \N__36195\,
            I => \N__36187\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__36190\,
            I => \N__36184\
        );

    \I__7476\ : Odrv4
    port map (
            O => \N__36187\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__7475\ : Odrv12
    port map (
            O => \N__36184\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__7474\ : InMux
    port map (
            O => \N__36179\,
            I => \bfn_16_10_0_\
        );

    \I__7473\ : CascadeMux
    port map (
            O => \N__36176\,
            I => \N__36173\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36170\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__36170\,
            I => \N__36165\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36169\,
            I => \N__36162\
        );

    \I__7469\ : InMux
    port map (
            O => \N__36168\,
            I => \N__36159\
        );

    \I__7468\ : Span4Mux_v
    port map (
            O => \N__36165\,
            I => \N__36154\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__36162\,
            I => \N__36154\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__36159\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__7465\ : Odrv4
    port map (
            O => \N__36154\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__7464\ : InMux
    port map (
            O => \N__36149\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__7463\ : InMux
    port map (
            O => \N__36146\,
            I => \N__36139\
        );

    \I__7462\ : InMux
    port map (
            O => \N__36145\,
            I => \N__36139\
        );

    \I__7461\ : InMux
    port map (
            O => \N__36144\,
            I => \N__36136\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__36139\,
            I => \N__36133\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__36136\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__7458\ : Odrv4
    port map (
            O => \N__36133\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__7457\ : InMux
    port map (
            O => \N__36128\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__7456\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36118\
        );

    \I__7455\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36118\
        );

    \I__7454\ : InMux
    port map (
            O => \N__36123\,
            I => \N__36115\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__36118\,
            I => \N__36112\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__36115\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__7451\ : Odrv4
    port map (
            O => \N__36112\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36107\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__7449\ : CascadeMux
    port map (
            O => \N__36104\,
            I => \N__36100\
        );

    \I__7448\ : InMux
    port map (
            O => \N__36103\,
            I => \N__36096\
        );

    \I__7447\ : InMux
    port map (
            O => \N__36100\,
            I => \N__36093\
        );

    \I__7446\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36090\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__36096\,
            I => \N__36085\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__36093\,
            I => \N__36085\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__36090\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__7442\ : Odrv4
    port map (
            O => \N__36085\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36080\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__7440\ : CascadeMux
    port map (
            O => \N__36077\,
            I => \N__36073\
        );

    \I__7439\ : InMux
    port map (
            O => \N__36076\,
            I => \N__36069\
        );

    \I__7438\ : InMux
    port map (
            O => \N__36073\,
            I => \N__36066\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36072\,
            I => \N__36063\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36069\,
            I => \N__36058\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__36066\,
            I => \N__36058\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__36063\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__7433\ : Odrv4
    port map (
            O => \N__36058\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__7432\ : InMux
    port map (
            O => \N__36053\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__7431\ : CascadeMux
    port map (
            O => \N__36050\,
            I => \N__36046\
        );

    \I__7430\ : CascadeMux
    port map (
            O => \N__36049\,
            I => \N__36043\
        );

    \I__7429\ : InMux
    port map (
            O => \N__36046\,
            I => \N__36037\
        );

    \I__7428\ : InMux
    port map (
            O => \N__36043\,
            I => \N__36037\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36042\,
            I => \N__36034\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__36037\,
            I => \N__36031\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__36034\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__36031\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__7423\ : InMux
    port map (
            O => \N__36026\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__7422\ : CascadeMux
    port map (
            O => \N__36023\,
            I => \N__36019\
        );

    \I__7421\ : CascadeMux
    port map (
            O => \N__36022\,
            I => \N__36016\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36019\,
            I => \N__36010\
        );

    \I__7419\ : InMux
    port map (
            O => \N__36016\,
            I => \N__36010\
        );

    \I__7418\ : InMux
    port map (
            O => \N__36015\,
            I => \N__36007\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__36010\,
            I => \N__36004\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__36007\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__7415\ : Odrv4
    port map (
            O => \N__36004\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__7414\ : InMux
    port map (
            O => \N__35999\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__7413\ : CascadeMux
    port map (
            O => \N__35996\,
            I => \N__35993\
        );

    \I__7412\ : InMux
    port map (
            O => \N__35993\,
            I => \N__35990\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__35990\,
            I => \N__35985\
        );

    \I__7410\ : InMux
    port map (
            O => \N__35989\,
            I => \N__35982\
        );

    \I__7409\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35979\
        );

    \I__7408\ : Span4Mux_v
    port map (
            O => \N__35985\,
            I => \N__35976\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__35982\,
            I => \N__35973\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__35979\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__7405\ : Odrv4
    port map (
            O => \N__35976\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__7404\ : Odrv4
    port map (
            O => \N__35973\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__7403\ : InMux
    port map (
            O => \N__35966\,
            I => \bfn_16_9_0_\
        );

    \I__7402\ : CascadeMux
    port map (
            O => \N__35963\,
            I => \N__35960\
        );

    \I__7401\ : InMux
    port map (
            O => \N__35960\,
            I => \N__35957\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__35957\,
            I => \N__35952\
        );

    \I__7399\ : InMux
    port map (
            O => \N__35956\,
            I => \N__35949\
        );

    \I__7398\ : InMux
    port map (
            O => \N__35955\,
            I => \N__35946\
        );

    \I__7397\ : Span4Mux_v
    port map (
            O => \N__35952\,
            I => \N__35941\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__35949\,
            I => \N__35941\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__35946\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__7394\ : Odrv4
    port map (
            O => \N__35941\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__7393\ : InMux
    port map (
            O => \N__35936\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__7392\ : CascadeMux
    port map (
            O => \N__35933\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\
        );

    \I__7391\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35927\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__35927\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\
        );

    \I__7389\ : CascadeMux
    port map (
            O => \N__35924\,
            I => \N__35920\
        );

    \I__7388\ : CascadeMux
    port map (
            O => \N__35923\,
            I => \N__35917\
        );

    \I__7387\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35914\
        );

    \I__7386\ : InMux
    port map (
            O => \N__35917\,
            I => \N__35910\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__35914\,
            I => \N__35907\
        );

    \I__7384\ : InMux
    port map (
            O => \N__35913\,
            I => \N__35904\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__35910\,
            I => \N__35897\
        );

    \I__7382\ : Span4Mux_v
    port map (
            O => \N__35907\,
            I => \N__35897\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__35904\,
            I => \N__35897\
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__35897\,
            I => \elapsed_time_ns_1_RNIAE2591_0_2\
        );

    \I__7379\ : CascadeMux
    port map (
            O => \N__35894\,
            I => \N__35891\
        );

    \I__7378\ : InMux
    port map (
            O => \N__35891\,
            I => \N__35887\
        );

    \I__7377\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35883\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__35887\,
            I => \N__35880\
        );

    \I__7375\ : InMux
    port map (
            O => \N__35886\,
            I => \N__35877\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__35883\,
            I => \N__35872\
        );

    \I__7373\ : Span4Mux_v
    port map (
            O => \N__35880\,
            I => \N__35872\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__35877\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__7371\ : Odrv4
    port map (
            O => \N__35872\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__7370\ : InMux
    port map (
            O => \N__35867\,
            I => \N__35864\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__35864\,
            I => \N__35861\
        );

    \I__7368\ : Span4Mux_h
    port map (
            O => \N__35861\,
            I => \N__35857\
        );

    \I__7367\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35854\
        );

    \I__7366\ : Odrv4
    port map (
            O => \N__35857\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__35854\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__7364\ : InMux
    port map (
            O => \N__35849\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__7363\ : InMux
    port map (
            O => \N__35846\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__7362\ : InMux
    port map (
            O => \N__35843\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__7361\ : InMux
    port map (
            O => \N__35840\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__7360\ : InMux
    port map (
            O => \N__35837\,
            I => \N__35834\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__35834\,
            I => \N__35831\
        );

    \I__7358\ : Span4Mux_h
    port map (
            O => \N__35831\,
            I => \N__35828\
        );

    \I__7357\ : Odrv4
    port map (
            O => \N__35828\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__7356\ : InMux
    port map (
            O => \N__35825\,
            I => \N__35822\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__35822\,
            I => \phase_controller_inst2.start_timer_hc_RNOZ0Z_0\
        );

    \I__7354\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35814\
        );

    \I__7353\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35811\
        );

    \I__7352\ : InMux
    port map (
            O => \N__35817\,
            I => \N__35807\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__35814\,
            I => \N__35804\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__35811\,
            I => \N__35801\
        );

    \I__7349\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35798\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__35807\,
            I => \N__35791\
        );

    \I__7347\ : Span12Mux_h
    port map (
            O => \N__35804\,
            I => \N__35791\
        );

    \I__7346\ : Span12Mux_s5_v
    port map (
            O => \N__35801\,
            I => \N__35791\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__35798\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7344\ : Odrv12
    port map (
            O => \N__35791\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7343\ : CEMux
    port map (
            O => \N__35786\,
            I => \N__35781\
        );

    \I__7342\ : CEMux
    port map (
            O => \N__35785\,
            I => \N__35778\
        );

    \I__7341\ : CEMux
    port map (
            O => \N__35784\,
            I => \N__35774\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__35781\,
            I => \N__35771\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__35778\,
            I => \N__35768\
        );

    \I__7338\ : CEMux
    port map (
            O => \N__35777\,
            I => \N__35765\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__35774\,
            I => \N__35762\
        );

    \I__7336\ : Span4Mux_v
    port map (
            O => \N__35771\,
            I => \N__35757\
        );

    \I__7335\ : Span4Mux_v
    port map (
            O => \N__35768\,
            I => \N__35757\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__35765\,
            I => \N__35754\
        );

    \I__7333\ : Span4Mux_v
    port map (
            O => \N__35762\,
            I => \N__35747\
        );

    \I__7332\ : Span4Mux_h
    port map (
            O => \N__35757\,
            I => \N__35747\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__35754\,
            I => \N__35747\
        );

    \I__7330\ : Odrv4
    port map (
            O => \N__35747\,
            I => \delay_measurement_inst.delay_tr_timer.N_435_i\
        );

    \I__7329\ : InMux
    port map (
            O => \N__35744\,
            I => \N__35738\
        );

    \I__7328\ : InMux
    port map (
            O => \N__35743\,
            I => \N__35733\
        );

    \I__7327\ : InMux
    port map (
            O => \N__35742\,
            I => \N__35733\
        );

    \I__7326\ : InMux
    port map (
            O => \N__35741\,
            I => \N__35730\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__35738\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__35733\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__35730\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7322\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35709\
        );

    \I__7321\ : InMux
    port map (
            O => \N__35722\,
            I => \N__35709\
        );

    \I__7320\ : InMux
    port map (
            O => \N__35721\,
            I => \N__35700\
        );

    \I__7319\ : InMux
    port map (
            O => \N__35720\,
            I => \N__35700\
        );

    \I__7318\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35700\
        );

    \I__7317\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35700\
        );

    \I__7316\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35687\
        );

    \I__7315\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35687\
        );

    \I__7314\ : InMux
    port map (
            O => \N__35715\,
            I => \N__35687\
        );

    \I__7313\ : InMux
    port map (
            O => \N__35714\,
            I => \N__35687\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__35709\,
            I => \N__35666\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__35700\,
            I => \N__35666\
        );

    \I__7310\ : InMux
    port map (
            O => \N__35699\,
            I => \N__35657\
        );

    \I__7309\ : InMux
    port map (
            O => \N__35698\,
            I => \N__35657\
        );

    \I__7308\ : InMux
    port map (
            O => \N__35697\,
            I => \N__35657\
        );

    \I__7307\ : InMux
    port map (
            O => \N__35696\,
            I => \N__35657\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__35687\,
            I => \N__35654\
        );

    \I__7305\ : InMux
    port map (
            O => \N__35686\,
            I => \N__35645\
        );

    \I__7304\ : InMux
    port map (
            O => \N__35685\,
            I => \N__35645\
        );

    \I__7303\ : InMux
    port map (
            O => \N__35684\,
            I => \N__35645\
        );

    \I__7302\ : InMux
    port map (
            O => \N__35683\,
            I => \N__35645\
        );

    \I__7301\ : InMux
    port map (
            O => \N__35682\,
            I => \N__35636\
        );

    \I__7300\ : InMux
    port map (
            O => \N__35681\,
            I => \N__35636\
        );

    \I__7299\ : InMux
    port map (
            O => \N__35680\,
            I => \N__35636\
        );

    \I__7298\ : InMux
    port map (
            O => \N__35679\,
            I => \N__35636\
        );

    \I__7297\ : InMux
    port map (
            O => \N__35678\,
            I => \N__35627\
        );

    \I__7296\ : InMux
    port map (
            O => \N__35677\,
            I => \N__35627\
        );

    \I__7295\ : InMux
    port map (
            O => \N__35676\,
            I => \N__35627\
        );

    \I__7294\ : InMux
    port map (
            O => \N__35675\,
            I => \N__35627\
        );

    \I__7293\ : InMux
    port map (
            O => \N__35674\,
            I => \N__35618\
        );

    \I__7292\ : InMux
    port map (
            O => \N__35673\,
            I => \N__35618\
        );

    \I__7291\ : InMux
    port map (
            O => \N__35672\,
            I => \N__35618\
        );

    \I__7290\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35618\
        );

    \I__7289\ : Span4Mux_h
    port map (
            O => \N__35666\,
            I => \N__35615\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__35657\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7287\ : Odrv4
    port map (
            O => \N__35654\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__35645\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__35636\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__35627\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__35618\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7282\ : Odrv4
    port map (
            O => \N__35615\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7281\ : InMux
    port map (
            O => \N__35600\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__7280\ : InMux
    port map (
            O => \N__35597\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__7279\ : InMux
    port map (
            O => \N__35594\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__7278\ : InMux
    port map (
            O => \N__35591\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__7277\ : InMux
    port map (
            O => \N__35588\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__7276\ : InMux
    port map (
            O => \N__35585\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__7275\ : InMux
    port map (
            O => \N__35582\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__7274\ : InMux
    port map (
            O => \N__35579\,
            I => \bfn_15_23_0_\
        );

    \I__7273\ : InMux
    port map (
            O => \N__35576\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__7272\ : CascadeMux
    port map (
            O => \N__35573\,
            I => \N__35569\
        );

    \I__7271\ : InMux
    port map (
            O => \N__35572\,
            I => \N__35565\
        );

    \I__7270\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35562\
        );

    \I__7269\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35559\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__35565\,
            I => \N__35556\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__35562\,
            I => \N__35551\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__35559\,
            I => \N__35551\
        );

    \I__7265\ : Span4Mux_v
    port map (
            O => \N__35556\,
            I => \N__35547\
        );

    \I__7264\ : Span4Mux_v
    port map (
            O => \N__35551\,
            I => \N__35544\
        );

    \I__7263\ : InMux
    port map (
            O => \N__35550\,
            I => \N__35541\
        );

    \I__7262\ : Odrv4
    port map (
            O => \N__35547\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__7261\ : Odrv4
    port map (
            O => \N__35544\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__35541\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__7259\ : InMux
    port map (
            O => \N__35534\,
            I => \bfn_15_21_0_\
        );

    \I__7258\ : InMux
    port map (
            O => \N__35531\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__7257\ : InMux
    port map (
            O => \N__35528\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__7256\ : InMux
    port map (
            O => \N__35525\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__7255\ : InMux
    port map (
            O => \N__35522\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__7254\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35516\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__35516\,
            I => \N__35512\
        );

    \I__7252\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35509\
        );

    \I__7251\ : Span4Mux_h
    port map (
            O => \N__35512\,
            I => \N__35503\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__35509\,
            I => \N__35503\
        );

    \I__7249\ : InMux
    port map (
            O => \N__35508\,
            I => \N__35500\
        );

    \I__7248\ : Span4Mux_v
    port map (
            O => \N__35503\,
            I => \N__35496\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__35500\,
            I => \N__35493\
        );

    \I__7246\ : InMux
    port map (
            O => \N__35499\,
            I => \N__35490\
        );

    \I__7245\ : Odrv4
    port map (
            O => \N__35496\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__7244\ : Odrv4
    port map (
            O => \N__35493\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__35490\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__7242\ : InMux
    port map (
            O => \N__35483\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__7241\ : InMux
    port map (
            O => \N__35480\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__7240\ : InMux
    port map (
            O => \N__35477\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__7239\ : InMux
    port map (
            O => \N__35474\,
            I => \N__35467\
        );

    \I__7238\ : InMux
    port map (
            O => \N__35473\,
            I => \N__35467\
        );

    \I__7237\ : CascadeMux
    port map (
            O => \N__35472\,
            I => \N__35464\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__35467\,
            I => \N__35461\
        );

    \I__7235\ : InMux
    port map (
            O => \N__35464\,
            I => \N__35458\
        );

    \I__7234\ : Span4Mux_h
    port map (
            O => \N__35461\,
            I => \N__35452\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__35458\,
            I => \N__35452\
        );

    \I__7232\ : InMux
    port map (
            O => \N__35457\,
            I => \N__35449\
        );

    \I__7231\ : Odrv4
    port map (
            O => \N__35452\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__35449\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__7229\ : InMux
    port map (
            O => \N__35444\,
            I => \bfn_15_22_0_\
        );

    \I__7228\ : CascadeMux
    port map (
            O => \N__35441\,
            I => \N__35438\
        );

    \I__7227\ : InMux
    port map (
            O => \N__35438\,
            I => \N__35431\
        );

    \I__7226\ : InMux
    port map (
            O => \N__35437\,
            I => \N__35431\
        );

    \I__7225\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35428\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__35431\,
            I => \N__35424\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__35428\,
            I => \N__35421\
        );

    \I__7222\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35418\
        );

    \I__7221\ : Span4Mux_v
    port map (
            O => \N__35424\,
            I => \N__35415\
        );

    \I__7220\ : Span4Mux_h
    port map (
            O => \N__35421\,
            I => \N__35412\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__35418\,
            I => \N__35409\
        );

    \I__7218\ : Odrv4
    port map (
            O => \N__35415\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__7217\ : Odrv4
    port map (
            O => \N__35412\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__7216\ : Odrv4
    port map (
            O => \N__35409\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__7215\ : InMux
    port map (
            O => \N__35402\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__7214\ : CascadeMux
    port map (
            O => \N__35399\,
            I => \N__35396\
        );

    \I__7213\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35392\
        );

    \I__7212\ : CascadeMux
    port map (
            O => \N__35395\,
            I => \N__35389\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__35392\,
            I => \N__35386\
        );

    \I__7210\ : InMux
    port map (
            O => \N__35389\,
            I => \N__35383\
        );

    \I__7209\ : Span4Mux_v
    port map (
            O => \N__35386\,
            I => \N__35376\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__35383\,
            I => \N__35376\
        );

    \I__7207\ : InMux
    port map (
            O => \N__35382\,
            I => \N__35373\
        );

    \I__7206\ : InMux
    port map (
            O => \N__35381\,
            I => \N__35370\
        );

    \I__7205\ : Span4Mux_h
    port map (
            O => \N__35376\,
            I => \N__35365\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__35373\,
            I => \N__35365\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__35370\,
            I => \N__35362\
        );

    \I__7202\ : Span4Mux_v
    port map (
            O => \N__35365\,
            I => \N__35359\
        );

    \I__7201\ : Span4Mux_h
    port map (
            O => \N__35362\,
            I => \N__35356\
        );

    \I__7200\ : Odrv4
    port map (
            O => \N__35359\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__7199\ : Odrv4
    port map (
            O => \N__35356\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__7198\ : InMux
    port map (
            O => \N__35351\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__7197\ : CascadeMux
    port map (
            O => \N__35348\,
            I => \N__35345\
        );

    \I__7196\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35341\
        );

    \I__7195\ : CascadeMux
    port map (
            O => \N__35344\,
            I => \N__35338\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__35341\,
            I => \N__35333\
        );

    \I__7193\ : InMux
    port map (
            O => \N__35338\,
            I => \N__35328\
        );

    \I__7192\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35328\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35336\,
            I => \N__35325\
        );

    \I__7190\ : Span4Mux_v
    port map (
            O => \N__35333\,
            I => \N__35320\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__35328\,
            I => \N__35320\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__35325\,
            I => \N__35317\
        );

    \I__7187\ : Span4Mux_v
    port map (
            O => \N__35320\,
            I => \N__35314\
        );

    \I__7186\ : Span4Mux_h
    port map (
            O => \N__35317\,
            I => \N__35311\
        );

    \I__7185\ : Odrv4
    port map (
            O => \N__35314\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__7184\ : Odrv4
    port map (
            O => \N__35311\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__7183\ : InMux
    port map (
            O => \N__35306\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__7182\ : InMux
    port map (
            O => \N__35303\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__7181\ : InMux
    port map (
            O => \N__35300\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__7180\ : InMux
    port map (
            O => \N__35297\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__7179\ : CascadeMux
    port map (
            O => \N__35294\,
            I => \N__35290\
        );

    \I__7178\ : InMux
    port map (
            O => \N__35293\,
            I => \N__35287\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35290\,
            I => \N__35284\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__35287\,
            I => \N__35279\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__35284\,
            I => \N__35279\
        );

    \I__7174\ : Span4Mux_v
    port map (
            O => \N__35279\,
            I => \N__35275\
        );

    \I__7173\ : InMux
    port map (
            O => \N__35278\,
            I => \N__35271\
        );

    \I__7172\ : Span4Mux_v
    port map (
            O => \N__35275\,
            I => \N__35268\
        );

    \I__7171\ : InMux
    port map (
            O => \N__35274\,
            I => \N__35265\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__35271\,
            I => \N__35262\
        );

    \I__7169\ : Odrv4
    port map (
            O => \N__35268\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__35265\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__7167\ : Odrv4
    port map (
            O => \N__35262\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35255\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__7165\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35249\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__35249\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__7163\ : InMux
    port map (
            O => \N__35246\,
            I => \N__35241\
        );

    \I__7162\ : InMux
    port map (
            O => \N__35245\,
            I => \N__35238\
        );

    \I__7161\ : CascadeMux
    port map (
            O => \N__35244\,
            I => \N__35235\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__35241\,
            I => \N__35232\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__35238\,
            I => \N__35229\
        );

    \I__7158\ : InMux
    port map (
            O => \N__35235\,
            I => \N__35226\
        );

    \I__7157\ : Odrv4
    port map (
            O => \N__35232\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__7156\ : Odrv12
    port map (
            O => \N__35229\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__35226\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35216\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__35216\,
            I => \N__35213\
        );

    \I__7152\ : Odrv4
    port map (
            O => \N__35213\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__7151\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35207\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35207\,
            I => \N__35204\
        );

    \I__7149\ : Odrv4
    port map (
            O => \N__35204\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__7148\ : CascadeMux
    port map (
            O => \N__35201\,
            I => \N__35197\
        );

    \I__7147\ : CascadeMux
    port map (
            O => \N__35200\,
            I => \N__35194\
        );

    \I__7146\ : InMux
    port map (
            O => \N__35197\,
            I => \N__35188\
        );

    \I__7145\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35188\
        );

    \I__7144\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35185\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__35188\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__35185\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35180\,
            I => \N__35177\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__35177\,
            I => \N__35174\
        );

    \I__7139\ : Odrv4
    port map (
            O => \N__35174\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__7138\ : InMux
    port map (
            O => \N__35171\,
            I => \N__35168\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__35168\,
            I => \N__35165\
        );

    \I__7136\ : Span4Mux_h
    port map (
            O => \N__35165\,
            I => \N__35162\
        );

    \I__7135\ : Odrv4
    port map (
            O => \N__35162\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__7134\ : InMux
    port map (
            O => \N__35159\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35156\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35153\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__7131\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35147\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35147\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__7129\ : CascadeMux
    port map (
            O => \N__35144\,
            I => \N__35141\
        );

    \I__7128\ : InMux
    port map (
            O => \N__35141\,
            I => \N__35138\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__35138\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__7126\ : InMux
    port map (
            O => \N__35135\,
            I => \N__35131\
        );

    \I__7125\ : InMux
    port map (
            O => \N__35134\,
            I => \N__35128\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__35131\,
            I => \N__35122\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__35128\,
            I => \N__35122\
        );

    \I__7122\ : InMux
    port map (
            O => \N__35127\,
            I => \N__35119\
        );

    \I__7121\ : Odrv12
    port map (
            O => \N__35122\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__35119\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__7119\ : InMux
    port map (
            O => \N__35114\,
            I => \N__35110\
        );

    \I__7118\ : InMux
    port map (
            O => \N__35113\,
            I => \N__35107\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__35110\,
            I => \N__35103\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__35107\,
            I => \N__35100\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35106\,
            I => \N__35097\
        );

    \I__7114\ : Odrv4
    port map (
            O => \N__35103\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__7113\ : Odrv4
    port map (
            O => \N__35100\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__35097\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__7111\ : CascadeMux
    port map (
            O => \N__35090\,
            I => \N__35087\
        );

    \I__7110\ : InMux
    port map (
            O => \N__35087\,
            I => \N__35084\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__35084\,
            I => \N__35081\
        );

    \I__7108\ : Span12Mux_v
    port map (
            O => \N__35081\,
            I => \N__35078\
        );

    \I__7107\ : Odrv12
    port map (
            O => \N__35078\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__7106\ : InMux
    port map (
            O => \N__35075\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35072\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__7104\ : CascadeMux
    port map (
            O => \N__35069\,
            I => \N__35066\
        );

    \I__7103\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35063\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__35063\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__7101\ : InMux
    port map (
            O => \N__35060\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__7100\ : InMux
    port map (
            O => \N__35057\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__7099\ : InMux
    port map (
            O => \N__35054\,
            I => \bfn_15_17_0_\
        );

    \I__7098\ : InMux
    port map (
            O => \N__35051\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__35048\,
            I => \N__35045\
        );

    \I__7096\ : InMux
    port map (
            O => \N__35045\,
            I => \N__35042\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__35042\,
            I => \N__35039\
        );

    \I__7094\ : Span4Mux_v
    port map (
            O => \N__35039\,
            I => \N__35036\
        );

    \I__7093\ : Odrv4
    port map (
            O => \N__35036\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__7092\ : InMux
    port map (
            O => \N__35033\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__7091\ : InMux
    port map (
            O => \N__35030\,
            I => \N__35027\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__35027\,
            I => \N__35024\
        );

    \I__7089\ : Span4Mux_h
    port map (
            O => \N__35024\,
            I => \N__35021\
        );

    \I__7088\ : Odrv4
    port map (
            O => \N__35021\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35018\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__7086\ : InMux
    port map (
            O => \N__35015\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__7085\ : CascadeMux
    port map (
            O => \N__35012\,
            I => \N__35009\
        );

    \I__7084\ : InMux
    port map (
            O => \N__35009\,
            I => \N__35006\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__35006\,
            I => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\
        );

    \I__7082\ : InMux
    port map (
            O => \N__35003\,
            I => \N__35000\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__35000\,
            I => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\
        );

    \I__7080\ : CascadeMux
    port map (
            O => \N__34997\,
            I => \N__34994\
        );

    \I__7079\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34991\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__34991\,
            I => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\
        );

    \I__7077\ : InMux
    port map (
            O => \N__34988\,
            I => \N__34985\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__34985\,
            I => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\
        );

    \I__7075\ : CascadeMux
    port map (
            O => \N__34982\,
            I => \N__34979\
        );

    \I__7074\ : InMux
    port map (
            O => \N__34979\,
            I => \N__34976\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__34976\,
            I => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\
        );

    \I__7072\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34970\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__34970\,
            I => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__34967\,
            I => \N__34964\
        );

    \I__7069\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34961\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__34961\,
            I => \N__34958\
        );

    \I__7067\ : Span4Mux_v
    port map (
            O => \N__34958\,
            I => \N__34955\
        );

    \I__7066\ : Odrv4
    port map (
            O => \N__34955\,
            I => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\
        );

    \I__7065\ : InMux
    port map (
            O => \N__34952\,
            I => \N__34949\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__34949\,
            I => \N__34946\
        );

    \I__7063\ : Span4Mux_h
    port map (
            O => \N__34946\,
            I => \N__34943\
        );

    \I__7062\ : Odrv4
    port map (
            O => \N__34943\,
            I => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\
        );

    \I__7061\ : InMux
    port map (
            O => \N__34940\,
            I => \N__34937\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__34937\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__7059\ : CascadeMux
    port map (
            O => \N__34934\,
            I => \N__34931\
        );

    \I__7058\ : InMux
    port map (
            O => \N__34931\,
            I => \N__34928\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__34928\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__7056\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34922\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__34922\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__7054\ : CascadeMux
    port map (
            O => \N__34919\,
            I => \N__34916\
        );

    \I__7053\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34913\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__34913\,
            I => \N__34910\
        );

    \I__7051\ : Span12Mux_v
    port map (
            O => \N__34910\,
            I => \N__34907\
        );

    \I__7050\ : Odrv12
    port map (
            O => \N__34907\,
            I => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\
        );

    \I__7049\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34901\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__34901\,
            I => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\
        );

    \I__7047\ : CascadeMux
    port map (
            O => \N__34898\,
            I => \N__34895\
        );

    \I__7046\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34892\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__34892\,
            I => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\
        );

    \I__7044\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34886\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__34886\,
            I => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\
        );

    \I__7042\ : CascadeMux
    port map (
            O => \N__34883\,
            I => \N__34880\
        );

    \I__7041\ : InMux
    port map (
            O => \N__34880\,
            I => \N__34877\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__34877\,
            I => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\
        );

    \I__7039\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34871\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__34871\,
            I => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\
        );

    \I__7037\ : InMux
    port map (
            O => \N__34868\,
            I => \N__34865\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__34865\,
            I => \N__34862\
        );

    \I__7035\ : Span4Mux_v
    port map (
            O => \N__34862\,
            I => \N__34859\
        );

    \I__7034\ : Odrv4
    port map (
            O => \N__34859\,
            I => \phase_controller_inst1.stoper_tr.un6_running_17\
        );

    \I__7033\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34852\
        );

    \I__7032\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34849\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__34852\,
            I => \N__34846\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__34849\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__34846\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7028\ : CascadeMux
    port map (
            O => \N__34841\,
            I => \N__34838\
        );

    \I__7027\ : InMux
    port map (
            O => \N__34838\,
            I => \N__34835\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__34835\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__7025\ : CascadeMux
    port map (
            O => \N__34832\,
            I => \N__34829\
        );

    \I__7024\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34826\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__34826\,
            I => \N__34823\
        );

    \I__7022\ : Odrv12
    port map (
            O => \N__34823\,
            I => \phase_controller_inst1.stoper_tr.un6_running_18\
        );

    \I__7021\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34816\
        );

    \I__7020\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34813\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__34816\,
            I => \N__34810\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__34813\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__7017\ : Odrv4
    port map (
            O => \N__34810\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__7016\ : InMux
    port map (
            O => \N__34805\,
            I => \N__34802\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__34802\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__7014\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34795\
        );

    \I__7013\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34792\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__34795\,
            I => \N__34789\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__34792\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__7010\ : Odrv4
    port map (
            O => \N__34789\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__7009\ : CascadeMux
    port map (
            O => \N__34784\,
            I => \N__34781\
        );

    \I__7008\ : InMux
    port map (
            O => \N__34781\,
            I => \N__34778\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__34778\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__7006\ : InMux
    port map (
            O => \N__34775\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_19\
        );

    \I__7005\ : InMux
    port map (
            O => \N__34772\,
            I => \N__34768\
        );

    \I__7004\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34764\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__34768\,
            I => \N__34761\
        );

    \I__7002\ : InMux
    port map (
            O => \N__34767\,
            I => \N__34758\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__34764\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__34761\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__34758\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO\
        );

    \I__6998\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34748\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__34748\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__6996\ : CascadeMux
    port map (
            O => \N__34745\,
            I => \N__34742\
        );

    \I__6995\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34739\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__34739\,
            I => \N__34736\
        );

    \I__6993\ : Span4Mux_h
    port map (
            O => \N__34736\,
            I => \N__34733\
        );

    \I__6992\ : Odrv4
    port map (
            O => \N__34733\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__34730\,
            I => \N__34727\
        );

    \I__6990\ : InMux
    port map (
            O => \N__34727\,
            I => \N__34724\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__34724\,
            I => \N__34721\
        );

    \I__6988\ : Odrv4
    port map (
            O => \N__34721\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__6987\ : InMux
    port map (
            O => \N__34718\,
            I => \N__34715\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__34715\,
            I => \N__34712\
        );

    \I__6985\ : Odrv12
    port map (
            O => \N__34712\,
            I => \phase_controller_inst1.stoper_tr.un6_running_10\
        );

    \I__6984\ : InMux
    port map (
            O => \N__34709\,
            I => \N__34705\
        );

    \I__6983\ : InMux
    port map (
            O => \N__34708\,
            I => \N__34702\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__34705\,
            I => \N__34699\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__34702\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__6980\ : Odrv4
    port map (
            O => \N__34699\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__6979\ : CascadeMux
    port map (
            O => \N__34694\,
            I => \N__34691\
        );

    \I__6978\ : InMux
    port map (
            O => \N__34691\,
            I => \N__34688\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__34688\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__6976\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34682\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__34682\,
            I => \N__34679\
        );

    \I__6974\ : Odrv4
    port map (
            O => \N__34679\,
            I => \phase_controller_inst1.stoper_tr.un6_running_11\
        );

    \I__6973\ : InMux
    port map (
            O => \N__34676\,
            I => \N__34672\
        );

    \I__6972\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34669\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__34672\,
            I => \N__34664\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__34669\,
            I => \N__34664\
        );

    \I__6969\ : Odrv4
    port map (
            O => \N__34664\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__6968\ : CascadeMux
    port map (
            O => \N__34661\,
            I => \N__34658\
        );

    \I__6967\ : InMux
    port map (
            O => \N__34658\,
            I => \N__34655\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__34655\,
            I => \N__34652\
        );

    \I__6965\ : Odrv4
    port map (
            O => \N__34652\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__6964\ : CascadeMux
    port map (
            O => \N__34649\,
            I => \N__34646\
        );

    \I__6963\ : InMux
    port map (
            O => \N__34646\,
            I => \N__34643\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__34643\,
            I => \N__34640\
        );

    \I__6961\ : Sp12to4
    port map (
            O => \N__34640\,
            I => \N__34637\
        );

    \I__6960\ : Odrv12
    port map (
            O => \N__34637\,
            I => \phase_controller_inst1.stoper_tr.un6_running_12\
        );

    \I__6959\ : InMux
    port map (
            O => \N__34634\,
            I => \N__34630\
        );

    \I__6958\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34627\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__34630\,
            I => \N__34622\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__34627\,
            I => \N__34622\
        );

    \I__6955\ : Odrv4
    port map (
            O => \N__34622\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__6954\ : InMux
    port map (
            O => \N__34619\,
            I => \N__34616\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__34616\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__6952\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34609\
        );

    \I__6951\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34606\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__34609\,
            I => \N__34603\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__34606\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__6948\ : Odrv4
    port map (
            O => \N__34603\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__6947\ : CascadeMux
    port map (
            O => \N__34598\,
            I => \N__34595\
        );

    \I__6946\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34592\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__34592\,
            I => \N__34589\
        );

    \I__6944\ : Odrv4
    port map (
            O => \N__34589\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__6943\ : InMux
    port map (
            O => \N__34586\,
            I => \N__34582\
        );

    \I__6942\ : InMux
    port map (
            O => \N__34585\,
            I => \N__34579\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__34582\,
            I => \N__34576\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__34579\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__6939\ : Odrv4
    port map (
            O => \N__34576\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__6938\ : CascadeMux
    port map (
            O => \N__34571\,
            I => \N__34568\
        );

    \I__6937\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34565\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__34565\,
            I => \N__34562\
        );

    \I__6935\ : Odrv4
    port map (
            O => \N__34562\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__6934\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34555\
        );

    \I__6933\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34552\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__34555\,
            I => \N__34549\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__34552\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__34549\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__6929\ : InMux
    port map (
            O => \N__34544\,
            I => \N__34541\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__34541\,
            I => \N__34538\
        );

    \I__6927\ : Span4Mux_v
    port map (
            O => \N__34538\,
            I => \N__34535\
        );

    \I__6926\ : Odrv4
    port map (
            O => \N__34535\,
            I => \phase_controller_inst1.stoper_tr.un6_running_15\
        );

    \I__6925\ : CascadeMux
    port map (
            O => \N__34532\,
            I => \N__34529\
        );

    \I__6924\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34526\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__34526\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__6922\ : InMux
    port map (
            O => \N__34523\,
            I => \N__34519\
        );

    \I__6921\ : InMux
    port map (
            O => \N__34522\,
            I => \N__34516\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__34519\,
            I => \N__34513\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__34516\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6918\ : Odrv4
    port map (
            O => \N__34513\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6917\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34505\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34502\
        );

    \I__6915\ : Span4Mux_v
    port map (
            O => \N__34502\,
            I => \N__34499\
        );

    \I__6914\ : Odrv4
    port map (
            O => \N__34499\,
            I => \phase_controller_inst1.stoper_tr.un6_running_16\
        );

    \I__6913\ : CascadeMux
    port map (
            O => \N__34496\,
            I => \N__34493\
        );

    \I__6912\ : InMux
    port map (
            O => \N__34493\,
            I => \N__34490\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__34490\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__6910\ : CascadeMux
    port map (
            O => \N__34487\,
            I => \N__34484\
        );

    \I__6909\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34481\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__34481\,
            I => \N__34478\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__34478\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__6906\ : InMux
    port map (
            O => \N__34475\,
            I => \N__34472\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__34472\,
            I => \N__34469\
        );

    \I__6904\ : Span4Mux_v
    port map (
            O => \N__34469\,
            I => \N__34466\
        );

    \I__6903\ : Odrv4
    port map (
            O => \N__34466\,
            I => \phase_controller_inst1.stoper_tr.un6_running_3\
        );

    \I__6902\ : InMux
    port map (
            O => \N__34463\,
            I => \N__34459\
        );

    \I__6901\ : InMux
    port map (
            O => \N__34462\,
            I => \N__34456\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__34459\,
            I => \N__34451\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__34456\,
            I => \N__34451\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__34451\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__6897\ : CascadeMux
    port map (
            O => \N__34448\,
            I => \N__34445\
        );

    \I__6896\ : InMux
    port map (
            O => \N__34445\,
            I => \N__34442\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34442\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__6894\ : InMux
    port map (
            O => \N__34439\,
            I => \N__34436\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__34436\,
            I => \N__34433\
        );

    \I__6892\ : Span4Mux_v
    port map (
            O => \N__34433\,
            I => \N__34430\
        );

    \I__6891\ : Odrv4
    port map (
            O => \N__34430\,
            I => \phase_controller_inst1.stoper_tr.un6_running_4\
        );

    \I__6890\ : InMux
    port map (
            O => \N__34427\,
            I => \N__34423\
        );

    \I__6889\ : InMux
    port map (
            O => \N__34426\,
            I => \N__34420\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__34423\,
            I => \N__34417\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__34420\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__6886\ : Odrv4
    port map (
            O => \N__34417\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__6885\ : CascadeMux
    port map (
            O => \N__34412\,
            I => \N__34409\
        );

    \I__6884\ : InMux
    port map (
            O => \N__34409\,
            I => \N__34406\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__34406\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__6882\ : InMux
    port map (
            O => \N__34403\,
            I => \N__34399\
        );

    \I__6881\ : InMux
    port map (
            O => \N__34402\,
            I => \N__34396\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__34399\,
            I => \N__34391\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__34396\,
            I => \N__34391\
        );

    \I__6878\ : Odrv4
    port map (
            O => \N__34391\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__6877\ : InMux
    port map (
            O => \N__34388\,
            I => \N__34385\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__34385\,
            I => \N__34382\
        );

    \I__6875\ : Span4Mux_v
    port map (
            O => \N__34382\,
            I => \N__34379\
        );

    \I__6874\ : Odrv4
    port map (
            O => \N__34379\,
            I => \phase_controller_inst1.stoper_tr.un6_running_5\
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__34376\,
            I => \N__34373\
        );

    \I__6872\ : InMux
    port map (
            O => \N__34373\,
            I => \N__34370\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__34370\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__6870\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34363\
        );

    \I__6869\ : InMux
    port map (
            O => \N__34366\,
            I => \N__34360\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__34363\,
            I => \N__34357\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__34360\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__6866\ : Odrv4
    port map (
            O => \N__34357\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__6865\ : InMux
    port map (
            O => \N__34352\,
            I => \N__34349\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__34349\,
            I => \N__34346\
        );

    \I__6863\ : Span4Mux_v
    port map (
            O => \N__34346\,
            I => \N__34343\
        );

    \I__6862\ : Odrv4
    port map (
            O => \N__34343\,
            I => \phase_controller_inst1.stoper_tr.un6_running_6\
        );

    \I__6861\ : CascadeMux
    port map (
            O => \N__34340\,
            I => \N__34337\
        );

    \I__6860\ : InMux
    port map (
            O => \N__34337\,
            I => \N__34334\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__34334\,
            I => \N__34331\
        );

    \I__6858\ : Odrv4
    port map (
            O => \N__34331\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__6857\ : InMux
    port map (
            O => \N__34328\,
            I => \N__34325\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__34325\,
            I => \N__34322\
        );

    \I__6855\ : Odrv4
    port map (
            O => \N__34322\,
            I => \phase_controller_inst1.stoper_tr.un6_running_7\
        );

    \I__6854\ : InMux
    port map (
            O => \N__34319\,
            I => \N__34315\
        );

    \I__6853\ : InMux
    port map (
            O => \N__34318\,
            I => \N__34312\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__34315\,
            I => \N__34309\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__34312\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__6850\ : Odrv12
    port map (
            O => \N__34309\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__6849\ : CascadeMux
    port map (
            O => \N__34304\,
            I => \N__34301\
        );

    \I__6848\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34298\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__34298\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__6846\ : InMux
    port map (
            O => \N__34295\,
            I => \N__34291\
        );

    \I__6845\ : InMux
    port map (
            O => \N__34294\,
            I => \N__34288\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__34291\,
            I => \N__34283\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__34288\,
            I => \N__34283\
        );

    \I__6842\ : Odrv4
    port map (
            O => \N__34283\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34280\,
            I => \N__34277\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34274\
        );

    \I__6839\ : Odrv12
    port map (
            O => \N__34274\,
            I => \phase_controller_inst1.stoper_tr.un6_running_8\
        );

    \I__6838\ : CascadeMux
    port map (
            O => \N__34271\,
            I => \N__34268\
        );

    \I__6837\ : InMux
    port map (
            O => \N__34268\,
            I => \N__34265\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__34265\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__6835\ : InMux
    port map (
            O => \N__34262\,
            I => \N__34259\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34259\,
            I => \N__34256\
        );

    \I__6833\ : Span4Mux_v
    port map (
            O => \N__34256\,
            I => \N__34253\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__34253\,
            I => \phase_controller_inst1.stoper_tr.un6_running_9\
        );

    \I__6831\ : InMux
    port map (
            O => \N__34250\,
            I => \N__34246\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34243\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__34246\,
            I => \N__34240\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__34243\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__34240\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__6826\ : CascadeMux
    port map (
            O => \N__34235\,
            I => \N__34232\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34232\,
            I => \N__34229\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__34229\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__6823\ : CascadeMux
    port map (
            O => \N__34226\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_\
        );

    \I__6822\ : InMux
    port map (
            O => \N__34223\,
            I => \N__34217\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34222\,
            I => \N__34214\
        );

    \I__6820\ : InMux
    port map (
            O => \N__34221\,
            I => \N__34211\
        );

    \I__6819\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34208\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__34217\,
            I => \phase_controller_inst1.stoper_tr.N_214\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__34214\,
            I => \phase_controller_inst1.stoper_tr.N_214\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__34211\,
            I => \phase_controller_inst1.stoper_tr.N_214\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__34208\,
            I => \phase_controller_inst1.stoper_tr.N_214\
        );

    \I__6814\ : CascadeMux
    port map (
            O => \N__34199\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34196\,
            I => \N__34193\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__34193\,
            I => \N__34187\
        );

    \I__6811\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34184\
        );

    \I__6810\ : CascadeMux
    port map (
            O => \N__34191\,
            I => \N__34181\
        );

    \I__6809\ : CascadeMux
    port map (
            O => \N__34190\,
            I => \N__34178\
        );

    \I__6808\ : Span4Mux_v
    port map (
            O => \N__34187\,
            I => \N__34174\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__34184\,
            I => \N__34171\
        );

    \I__6806\ : InMux
    port map (
            O => \N__34181\,
            I => \N__34166\
        );

    \I__6805\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34163\
        );

    \I__6804\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34160\
        );

    \I__6803\ : Sp12to4
    port map (
            O => \N__34174\,
            I => \N__34157\
        );

    \I__6802\ : Span4Mux_v
    port map (
            O => \N__34171\,
            I => \N__34154\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34170\,
            I => \N__34149\
        );

    \I__6800\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34149\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__34166\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__34163\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__34160\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__6796\ : Odrv12
    port map (
            O => \N__34157\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__6795\ : Odrv4
    port map (
            O => \N__34154\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34149\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__6793\ : CascadeMux
    port map (
            O => \N__34136\,
            I => \phase_controller_inst1.stoper_tr.N_241_cascade_\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34133\,
            I => \N__34130\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34130\,
            I => \N__34127\
        );

    \I__6790\ : Span4Mux_v
    port map (
            O => \N__34127\,
            I => \N__34124\
        );

    \I__6789\ : Odrv4
    port map (
            O => \N__34124\,
            I => \phase_controller_inst1.stoper_tr.un6_running_1\
        );

    \I__6788\ : CascadeMux
    port map (
            O => \N__34121\,
            I => \N__34117\
        );

    \I__6787\ : CascadeMux
    port map (
            O => \N__34120\,
            I => \N__34114\
        );

    \I__6786\ : InMux
    port map (
            O => \N__34117\,
            I => \N__34111\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34107\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__34111\,
            I => \N__34104\
        );

    \I__6783\ : InMux
    port map (
            O => \N__34110\,
            I => \N__34101\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__34107\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6781\ : Odrv4
    port map (
            O => \N__34104\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__34101\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6779\ : CascadeMux
    port map (
            O => \N__34094\,
            I => \N__34091\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34091\,
            I => \N__34088\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__34088\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__6776\ : InMux
    port map (
            O => \N__34085\,
            I => \N__34082\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__34082\,
            I => \N__34079\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__34079\,
            I => \N__34076\
        );

    \I__6773\ : Odrv4
    port map (
            O => \N__34076\,
            I => \phase_controller_inst1.stoper_tr.un6_running_2\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34069\
        );

    \I__6771\ : InMux
    port map (
            O => \N__34072\,
            I => \N__34066\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__34069\,
            I => \N__34063\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__34066\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__34063\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34058\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34055\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34052\,
            I => \N__34046\
        );

    \I__6764\ : InMux
    port map (
            O => \N__34051\,
            I => \N__34043\
        );

    \I__6763\ : InMux
    port map (
            O => \N__34050\,
            I => \N__34040\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34049\,
            I => \N__34037\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__34046\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__34043\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__34040\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__34037\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34028\,
            I => \N__34022\
        );

    \I__6756\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34019\
        );

    \I__6755\ : InMux
    port map (
            O => \N__34026\,
            I => \N__34014\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34025\,
            I => \N__34014\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__34022\,
            I => \elapsed_time_ns_1_RNIHI4DM1_0_18\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__34019\,
            I => \elapsed_time_ns_1_RNIHI4DM1_0_18\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__34014\,
            I => \elapsed_time_ns_1_RNIHI4DM1_0_18\
        );

    \I__6750\ : InMux
    port map (
            O => \N__34007\,
            I => \N__34004\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__34004\,
            I => \N__33988\
        );

    \I__6748\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33983\
        );

    \I__6747\ : InMux
    port map (
            O => \N__34002\,
            I => \N__33983\
        );

    \I__6746\ : InMux
    port map (
            O => \N__34001\,
            I => \N__33980\
        );

    \I__6745\ : InMux
    port map (
            O => \N__34000\,
            I => \N__33973\
        );

    \I__6744\ : InMux
    port map (
            O => \N__33999\,
            I => \N__33973\
        );

    \I__6743\ : InMux
    port map (
            O => \N__33998\,
            I => \N__33973\
        );

    \I__6742\ : InMux
    port map (
            O => \N__33997\,
            I => \N__33966\
        );

    \I__6741\ : InMux
    port map (
            O => \N__33996\,
            I => \N__33966\
        );

    \I__6740\ : InMux
    port map (
            O => \N__33995\,
            I => \N__33966\
        );

    \I__6739\ : InMux
    port map (
            O => \N__33994\,
            I => \N__33957\
        );

    \I__6738\ : InMux
    port map (
            O => \N__33993\,
            I => \N__33957\
        );

    \I__6737\ : InMux
    port map (
            O => \N__33992\,
            I => \N__33957\
        );

    \I__6736\ : InMux
    port map (
            O => \N__33991\,
            I => \N__33957\
        );

    \I__6735\ : Span4Mux_h
    port map (
            O => \N__33988\,
            I => \N__33954\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__33983\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__33980\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__33973\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__33966\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__33957\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__6729\ : Odrv4
    port map (
            O => \N__33954\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__6728\ : InMux
    port map (
            O => \N__33941\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__6727\ : InMux
    port map (
            O => \N__33938\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__6726\ : InMux
    port map (
            O => \N__33935\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__6725\ : InMux
    port map (
            O => \N__33932\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__6724\ : InMux
    port map (
            O => \N__33929\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__6723\ : InMux
    port map (
            O => \N__33926\,
            I => \bfn_15_8_0_\
        );

    \I__6722\ : InMux
    port map (
            O => \N__33923\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__6721\ : InMux
    port map (
            O => \N__33920\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__6720\ : InMux
    port map (
            O => \N__33917\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__6719\ : InMux
    port map (
            O => \N__33914\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__6718\ : InMux
    port map (
            O => \N__33911\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__6717\ : InMux
    port map (
            O => \N__33908\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__6716\ : InMux
    port map (
            O => \N__33905\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__6715\ : InMux
    port map (
            O => \N__33902\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__6714\ : InMux
    port map (
            O => \N__33899\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__6713\ : InMux
    port map (
            O => \N__33896\,
            I => \bfn_15_7_0_\
        );

    \I__6712\ : InMux
    port map (
            O => \N__33893\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__6711\ : InMux
    port map (
            O => \N__33890\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__6710\ : InMux
    port map (
            O => \N__33887\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__6709\ : InMux
    port map (
            O => \N__33884\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__6708\ : InMux
    port map (
            O => \N__33881\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__6707\ : InMux
    port map (
            O => \N__33878\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__6706\ : InMux
    port map (
            O => \N__33875\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33872\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__6704\ : InMux
    port map (
            O => \N__33869\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__6703\ : InMux
    port map (
            O => \N__33866\,
            I => \bfn_15_6_0_\
        );

    \I__6702\ : InMux
    port map (
            O => \N__33863\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__6701\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33857\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__33857\,
            I => \N__33854\
        );

    \I__6699\ : Odrv4
    port map (
            O => \N__33854\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__6698\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33848\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__33848\,
            I => \N__33845\
        );

    \I__6696\ : Odrv4
    port map (
            O => \N__33845\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__6695\ : InMux
    port map (
            O => \N__33842\,
            I => \N__33839\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__33839\,
            I => \N__33836\
        );

    \I__6693\ : Odrv4
    port map (
            O => \N__33836\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__6692\ : InMux
    port map (
            O => \N__33833\,
            I => \N__33830\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__33830\,
            I => \N__33827\
        );

    \I__6690\ : Odrv4
    port map (
            O => \N__33827\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__6689\ : InMux
    port map (
            O => \N__33824\,
            I => \N__33820\
        );

    \I__6688\ : CascadeMux
    port map (
            O => \N__33823\,
            I => \N__33817\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__33820\,
            I => \N__33813\
        );

    \I__6686\ : InMux
    port map (
            O => \N__33817\,
            I => \N__33810\
        );

    \I__6685\ : InMux
    port map (
            O => \N__33816\,
            I => \N__33807\
        );

    \I__6684\ : Odrv4
    port map (
            O => \N__33813\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__33810\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__33807\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__6681\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33797\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__33797\,
            I => \N__33793\
        );

    \I__6679\ : InMux
    port map (
            O => \N__33796\,
            I => \N__33790\
        );

    \I__6678\ : Span4Mux_v
    port map (
            O => \N__33793\,
            I => \N__33787\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__33790\,
            I => \N__33784\
        );

    \I__6676\ : Span4Mux_h
    port map (
            O => \N__33787\,
            I => \N__33781\
        );

    \I__6675\ : Span4Mux_h
    port map (
            O => \N__33784\,
            I => \N__33778\
        );

    \I__6674\ : Odrv4
    port map (
            O => \N__33781\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__6673\ : Odrv4
    port map (
            O => \N__33778\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__6672\ : CEMux
    port map (
            O => \N__33773\,
            I => \N__33755\
        );

    \I__6671\ : CEMux
    port map (
            O => \N__33772\,
            I => \N__33755\
        );

    \I__6670\ : CEMux
    port map (
            O => \N__33771\,
            I => \N__33755\
        );

    \I__6669\ : CEMux
    port map (
            O => \N__33770\,
            I => \N__33755\
        );

    \I__6668\ : CEMux
    port map (
            O => \N__33769\,
            I => \N__33755\
        );

    \I__6667\ : CEMux
    port map (
            O => \N__33768\,
            I => \N__33755\
        );

    \I__6666\ : GlobalMux
    port map (
            O => \N__33755\,
            I => \N__33752\
        );

    \I__6665\ : gio2CtrlBuf
    port map (
            O => \N__33752\,
            I => \delay_measurement_inst.delay_hc_timer.N_432_i_g\
        );

    \I__6664\ : CascadeMux
    port map (
            O => \N__33749\,
            I => \N__33743\
        );

    \I__6663\ : InMux
    port map (
            O => \N__33748\,
            I => \N__33740\
        );

    \I__6662\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33735\
        );

    \I__6661\ : InMux
    port map (
            O => \N__33746\,
            I => \N__33735\
        );

    \I__6660\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33732\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__33740\,
            I => \N__33727\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__33735\,
            I => \N__33727\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__33732\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6656\ : Odrv4
    port map (
            O => \N__33727\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6655\ : InMux
    port map (
            O => \N__33722\,
            I => \N__33719\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__33719\,
            I => \N__33716\
        );

    \I__6653\ : Span4Mux_h
    port map (
            O => \N__33716\,
            I => \N__33711\
        );

    \I__6652\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33708\
        );

    \I__6651\ : InMux
    port map (
            O => \N__33714\,
            I => \N__33705\
        );

    \I__6650\ : Span4Mux_v
    port map (
            O => \N__33711\,
            I => \N__33702\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__33708\,
            I => \N__33699\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__33705\,
            I => \N__33696\
        );

    \I__6647\ : Sp12to4
    port map (
            O => \N__33702\,
            I => \N__33689\
        );

    \I__6646\ : Sp12to4
    port map (
            O => \N__33699\,
            I => \N__33689\
        );

    \I__6645\ : Span12Mux_s9_v
    port map (
            O => \N__33696\,
            I => \N__33689\
        );

    \I__6644\ : Span12Mux_v
    port map (
            O => \N__33689\,
            I => \N__33686\
        );

    \I__6643\ : Odrv12
    port map (
            O => \N__33686\,
            I => \il_max_comp2_D2\
        );

    \I__6642\ : InMux
    port map (
            O => \N__33683\,
            I => \N__33680\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__33680\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__6640\ : IoInMux
    port map (
            O => \N__33677\,
            I => \N__33674\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__33674\,
            I => \N__33671\
        );

    \I__6638\ : Span4Mux_s3_v
    port map (
            O => \N__33671\,
            I => \N__33668\
        );

    \I__6637\ : Odrv4
    port map (
            O => \N__33668\,
            I => \delay_measurement_inst.delay_tr_timer.N_434_i\
        );

    \I__6636\ : InMux
    port map (
            O => \N__33665\,
            I => \bfn_15_5_0_\
        );

    \I__6635\ : InMux
    port map (
            O => \N__33662\,
            I => \N__33659\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__33659\,
            I => \N__33656\
        );

    \I__6633\ : Odrv4
    port map (
            O => \N__33656\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__6632\ : InMux
    port map (
            O => \N__33653\,
            I => \N__33650\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__33650\,
            I => \N__33647\
        );

    \I__6630\ : Span4Mux_h
    port map (
            O => \N__33647\,
            I => \N__33644\
        );

    \I__6629\ : Odrv4
    port map (
            O => \N__33644\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__6628\ : InMux
    port map (
            O => \N__33641\,
            I => \N__33638\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__33638\,
            I => \N__33635\
        );

    \I__6626\ : Odrv12
    port map (
            O => \N__33635\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__6625\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33629\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__33629\,
            I => \N__33626\
        );

    \I__6623\ : Odrv12
    port map (
            O => \N__33626\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__6622\ : InMux
    port map (
            O => \N__33623\,
            I => \N__33620\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__33620\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__6620\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33614\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__33614\,
            I => \N__33611\
        );

    \I__6618\ : Odrv4
    port map (
            O => \N__33611\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__6617\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33605\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__33605\,
            I => \N__33602\
        );

    \I__6615\ : Odrv12
    port map (
            O => \N__33602\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__6614\ : InMux
    port map (
            O => \N__33599\,
            I => \N__33596\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__33596\,
            I => \N__33593\
        );

    \I__6612\ : Odrv12
    port map (
            O => \N__33593\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__6611\ : InMux
    port map (
            O => \N__33590\,
            I => \N__33587\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__33587\,
            I => \N__33584\
        );

    \I__6609\ : Odrv12
    port map (
            O => \N__33584\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__6608\ : InMux
    port map (
            O => \N__33581\,
            I => \bfn_14_20_0_\
        );

    \I__6607\ : InMux
    port map (
            O => \N__33578\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__6606\ : InMux
    port map (
            O => \N__33575\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__6605\ : InMux
    port map (
            O => \N__33572\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__6604\ : InMux
    port map (
            O => \N__33569\,
            I => \N__33566\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__33566\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__6602\ : InMux
    port map (
            O => \N__33563\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33560\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__6600\ : CascadeMux
    port map (
            O => \N__33557\,
            I => \N__33554\
        );

    \I__6599\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33548\
        );

    \I__6598\ : InMux
    port map (
            O => \N__33553\,
            I => \N__33548\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__33548\,
            I => \N__33545\
        );

    \I__6596\ : Odrv4
    port map (
            O => \N__33545\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__6595\ : InMux
    port map (
            O => \N__33542\,
            I => \N__33539\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__33539\,
            I => \N__33536\
        );

    \I__6593\ : Odrv12
    port map (
            O => \N__33536\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__6592\ : InMux
    port map (
            O => \N__33533\,
            I => \N__33530\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__33530\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__6590\ : InMux
    port map (
            O => \N__33527\,
            I => \N__33524\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__33524\,
            I => \N__33521\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__33521\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__6587\ : InMux
    port map (
            O => \N__33518\,
            I => \N__33515\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__33515\,
            I => \N__33512\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__33512\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__6584\ : InMux
    port map (
            O => \N__33509\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__6583\ : InMux
    port map (
            O => \N__33506\,
            I => \bfn_14_19_0_\
        );

    \I__6582\ : InMux
    port map (
            O => \N__33503\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__6581\ : InMux
    port map (
            O => \N__33500\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__6580\ : InMux
    port map (
            O => \N__33497\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__6579\ : InMux
    port map (
            O => \N__33494\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__6578\ : InMux
    port map (
            O => \N__33491\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__6577\ : InMux
    port map (
            O => \N__33488\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__6576\ : InMux
    port map (
            O => \N__33485\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__6575\ : InMux
    port map (
            O => \N__33482\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__6574\ : InMux
    port map (
            O => \N__33479\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33473\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__33473\,
            I => \N__33470\
        );

    \I__6571\ : Span4Mux_v
    port map (
            O => \N__33470\,
            I => \N__33467\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__33467\,
            I => \N__33464\
        );

    \I__6569\ : Odrv4
    port map (
            O => \N__33464\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__6568\ : InMux
    port map (
            O => \N__33461\,
            I => \bfn_14_18_0_\
        );

    \I__6567\ : InMux
    port map (
            O => \N__33458\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__6566\ : InMux
    port map (
            O => \N__33455\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__6565\ : InMux
    port map (
            O => \N__33452\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__6564\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33446\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__33446\,
            I => \N__33443\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__33443\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__6561\ : InMux
    port map (
            O => \N__33440\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__6560\ : InMux
    port map (
            O => \N__33437\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__6559\ : InMux
    port map (
            O => \N__33434\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__6558\ : InMux
    port map (
            O => \N__33431\,
            I => \N__33428\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__33428\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__6556\ : CascadeMux
    port map (
            O => \N__33425\,
            I => \N__33422\
        );

    \I__6555\ : InMux
    port map (
            O => \N__33422\,
            I => \N__33418\
        );

    \I__6554\ : InMux
    port map (
            O => \N__33421\,
            I => \N__33414\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__33418\,
            I => \N__33411\
        );

    \I__6552\ : CascadeMux
    port map (
            O => \N__33417\,
            I => \N__33407\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__33414\,
            I => \N__33404\
        );

    \I__6550\ : Span4Mux_v
    port map (
            O => \N__33411\,
            I => \N__33401\
        );

    \I__6549\ : InMux
    port map (
            O => \N__33410\,
            I => \N__33398\
        );

    \I__6548\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33395\
        );

    \I__6547\ : Odrv4
    port map (
            O => \N__33404\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__6546\ : Odrv4
    port map (
            O => \N__33401\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__33398\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__33395\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__6543\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33377\
        );

    \I__6542\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33377\
        );

    \I__6541\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33377\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__33377\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__6539\ : InMux
    port map (
            O => \N__33374\,
            I => \N__33368\
        );

    \I__6538\ : InMux
    port map (
            O => \N__33373\,
            I => \N__33368\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__33368\,
            I => \N__33364\
        );

    \I__6536\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33361\
        );

    \I__6535\ : Odrv4
    port map (
            O => \N__33364\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__33361\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33356\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__6532\ : InMux
    port map (
            O => \N__33353\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__6531\ : InMux
    port map (
            O => \N__33350\,
            I => \N__33347\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__33347\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__6529\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33341\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__33341\,
            I => \N__33336\
        );

    \I__6527\ : InMux
    port map (
            O => \N__33340\,
            I => \N__33333\
        );

    \I__6526\ : InMux
    port map (
            O => \N__33339\,
            I => \N__33330\
        );

    \I__6525\ : Odrv4
    port map (
            O => \N__33336\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__33333\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__33330\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__6522\ : InMux
    port map (
            O => \N__33323\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__6521\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33317\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__33317\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__6519\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33311\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__33311\,
            I => \N__33306\
        );

    \I__6517\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33301\
        );

    \I__6516\ : InMux
    port map (
            O => \N__33309\,
            I => \N__33301\
        );

    \I__6515\ : Odrv4
    port map (
            O => \N__33306\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__33301\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__6513\ : InMux
    port map (
            O => \N__33296\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__6512\ : InMux
    port map (
            O => \N__33293\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__6511\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33287\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__33287\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__6509\ : CascadeMux
    port map (
            O => \N__33284\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__6508\ : InMux
    port map (
            O => \N__33281\,
            I => \N__33278\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__33278\,
            I => \N__33273\
        );

    \I__6506\ : InMux
    port map (
            O => \N__33277\,
            I => \N__33270\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33276\,
            I => \N__33267\
        );

    \I__6504\ : Span4Mux_v
    port map (
            O => \N__33273\,
            I => \N__33264\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__33270\,
            I => \N__33258\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__33267\,
            I => \N__33258\
        );

    \I__6501\ : Span4Mux_h
    port map (
            O => \N__33264\,
            I => \N__33255\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33263\,
            I => \N__33252\
        );

    \I__6499\ : Odrv4
    port map (
            O => \N__33258\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6498\ : Odrv4
    port map (
            O => \N__33255\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__33252\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6496\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33241\
        );

    \I__6495\ : InMux
    port map (
            O => \N__33244\,
            I => \N__33238\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33235\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33229\
        );

    \I__6492\ : Span4Mux_v
    port map (
            O => \N__33235\,
            I => \N__33226\
        );

    \I__6491\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33219\
        );

    \I__6490\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33219\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33219\
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__33229\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__33226\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__33219\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6485\ : CascadeMux
    port map (
            O => \N__33212\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__6484\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33206\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__33206\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__6482\ : CascadeMux
    port map (
            O => \N__33203\,
            I => \N__33200\
        );

    \I__6481\ : InMux
    port map (
            O => \N__33200\,
            I => \N__33194\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33199\,
            I => \N__33191\
        );

    \I__6479\ : InMux
    port map (
            O => \N__33198\,
            I => \N__33186\
        );

    \I__6478\ : InMux
    port map (
            O => \N__33197\,
            I => \N__33186\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__33194\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__33191\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__33186\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6474\ : InMux
    port map (
            O => \N__33179\,
            I => \N__33175\
        );

    \I__6473\ : InMux
    port map (
            O => \N__33178\,
            I => \N__33172\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__33175\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33172\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__33167\,
            I => \N__33164\
        );

    \I__6469\ : InMux
    port map (
            O => \N__33164\,
            I => \N__33161\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__33161\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6NZ0Z32\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33158\,
            I => \N__33155\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__33155\,
            I => \N__33152\
        );

    \I__6465\ : Span4Mux_h
    port map (
            O => \N__33152\,
            I => \N__33149\
        );

    \I__6464\ : Span4Mux_h
    port map (
            O => \N__33149\,
            I => \N__33146\
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__33146\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__6462\ : InMux
    port map (
            O => \N__33143\,
            I => \N__33140\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__33140\,
            I => \N__33137\
        );

    \I__6460\ : Span4Mux_v
    port map (
            O => \N__33137\,
            I => \N__33122\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33117\
        );

    \I__6458\ : InMux
    port map (
            O => \N__33135\,
            I => \N__33117\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__33134\,
            I => \N__33113\
        );

    \I__6456\ : CascadeMux
    port map (
            O => \N__33133\,
            I => \N__33106\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__33132\,
            I => \N__33100\
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__33131\,
            I => \N__33097\
        );

    \I__6453\ : CascadeMux
    port map (
            O => \N__33130\,
            I => \N__33094\
        );

    \I__6452\ : CascadeMux
    port map (
            O => \N__33129\,
            I => \N__33091\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__33128\,
            I => \N__33085\
        );

    \I__6450\ : CascadeMux
    port map (
            O => \N__33127\,
            I => \N__33081\
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__33126\,
            I => \N__33077\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__33125\,
            I => \N__33070\
        );

    \I__6447\ : Span4Mux_h
    port map (
            O => \N__33122\,
            I => \N__33060\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__33060\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33057\
        );

    \I__6444\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33054\
        );

    \I__6443\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33051\
        );

    \I__6442\ : InMux
    port map (
            O => \N__33111\,
            I => \N__33043\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33030\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33109\,
            I => \N__33030\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33106\,
            I => \N__33030\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33105\,
            I => \N__33030\
        );

    \I__6437\ : InMux
    port map (
            O => \N__33104\,
            I => \N__33030\
        );

    \I__6436\ : InMux
    port map (
            O => \N__33103\,
            I => \N__33030\
        );

    \I__6435\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33027\
        );

    \I__6434\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33024\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33094\,
            I => \N__33011\
        );

    \I__6432\ : InMux
    port map (
            O => \N__33091\,
            I => \N__33011\
        );

    \I__6431\ : InMux
    port map (
            O => \N__33090\,
            I => \N__33011\
        );

    \I__6430\ : InMux
    port map (
            O => \N__33089\,
            I => \N__33011\
        );

    \I__6429\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33011\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33011\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33084\,
            I => \N__33008\
        );

    \I__6426\ : InMux
    port map (
            O => \N__33081\,
            I => \N__32993\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33080\,
            I => \N__32993\
        );

    \I__6424\ : InMux
    port map (
            O => \N__33077\,
            I => \N__32993\
        );

    \I__6423\ : InMux
    port map (
            O => \N__33076\,
            I => \N__32993\
        );

    \I__6422\ : InMux
    port map (
            O => \N__33075\,
            I => \N__32993\
        );

    \I__6421\ : InMux
    port map (
            O => \N__33074\,
            I => \N__32993\
        );

    \I__6420\ : InMux
    port map (
            O => \N__33073\,
            I => \N__32993\
        );

    \I__6419\ : InMux
    port map (
            O => \N__33070\,
            I => \N__32986\
        );

    \I__6418\ : InMux
    port map (
            O => \N__33069\,
            I => \N__32986\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33068\,
            I => \N__32986\
        );

    \I__6416\ : CascadeMux
    port map (
            O => \N__33067\,
            I => \N__32983\
        );

    \I__6415\ : CascadeMux
    port map (
            O => \N__33066\,
            I => \N__32979\
        );

    \I__6414\ : CascadeMux
    port map (
            O => \N__33065\,
            I => \N__32975\
        );

    \I__6413\ : Span4Mux_v
    port map (
            O => \N__33060\,
            I => \N__32965\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__33057\,
            I => \N__32965\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__33054\,
            I => \N__32965\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__33051\,
            I => \N__32965\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33050\,
            I => \N__32960\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33049\,
            I => \N__32960\
        );

    \I__6407\ : InMux
    port map (
            O => \N__33048\,
            I => \N__32957\
        );

    \I__6406\ : InMux
    port map (
            O => \N__33047\,
            I => \N__32954\
        );

    \I__6405\ : InMux
    port map (
            O => \N__33046\,
            I => \N__32951\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__33043\,
            I => \N__32938\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__33030\,
            I => \N__32938\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__33027\,
            I => \N__32927\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__33024\,
            I => \N__32927\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__33011\,
            I => \N__32927\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__33008\,
            I => \N__32927\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__32993\,
            I => \N__32927\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__32986\,
            I => \N__32924\
        );

    \I__6396\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32911\
        );

    \I__6395\ : InMux
    port map (
            O => \N__32982\,
            I => \N__32911\
        );

    \I__6394\ : InMux
    port map (
            O => \N__32979\,
            I => \N__32911\
        );

    \I__6393\ : InMux
    port map (
            O => \N__32978\,
            I => \N__32911\
        );

    \I__6392\ : InMux
    port map (
            O => \N__32975\,
            I => \N__32911\
        );

    \I__6391\ : InMux
    port map (
            O => \N__32974\,
            I => \N__32911\
        );

    \I__6390\ : Span4Mux_v
    port map (
            O => \N__32965\,
            I => \N__32904\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__32960\,
            I => \N__32904\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__32957\,
            I => \N__32904\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__32954\,
            I => \N__32899\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__32951\,
            I => \N__32899\
        );

    \I__6385\ : InMux
    port map (
            O => \N__32950\,
            I => \N__32882\
        );

    \I__6384\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32882\
        );

    \I__6383\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32882\
        );

    \I__6382\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32882\
        );

    \I__6381\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32882\
        );

    \I__6380\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32882\
        );

    \I__6379\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32882\
        );

    \I__6378\ : InMux
    port map (
            O => \N__32943\,
            I => \N__32882\
        );

    \I__6377\ : Span4Mux_v
    port map (
            O => \N__32938\,
            I => \N__32877\
        );

    \I__6376\ : Span4Mux_v
    port map (
            O => \N__32927\,
            I => \N__32877\
        );

    \I__6375\ : Span12Mux_v
    port map (
            O => \N__32924\,
            I => \N__32872\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__32911\,
            I => \N__32872\
        );

    \I__6373\ : Span4Mux_h
    port map (
            O => \N__32904\,
            I => \N__32869\
        );

    \I__6372\ : Odrv12
    port map (
            O => \N__32899\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__32882\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6370\ : Odrv4
    port map (
            O => \N__32877\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6369\ : Odrv12
    port map (
            O => \N__32872\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6368\ : Odrv4
    port map (
            O => \N__32869\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6367\ : CascadeMux
    port map (
            O => \N__32858\,
            I => \N__32854\
        );

    \I__6366\ : CascadeMux
    port map (
            O => \N__32857\,
            I => \N__32850\
        );

    \I__6365\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32843\
        );

    \I__6364\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32843\
        );

    \I__6363\ : InMux
    port map (
            O => \N__32850\,
            I => \N__32843\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__32843\,
            I => \N__32840\
        );

    \I__6361\ : Span4Mux_v
    port map (
            O => \N__32840\,
            I => \N__32837\
        );

    \I__6360\ : Odrv4
    port map (
            O => \N__32837\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_0_12\
        );

    \I__6359\ : CascadeMux
    port map (
            O => \N__32834\,
            I => \elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_\
        );

    \I__6358\ : CascadeMux
    port map (
            O => \N__32831\,
            I => \N__32827\
        );

    \I__6357\ : CascadeMux
    port map (
            O => \N__32830\,
            I => \N__32824\
        );

    \I__6356\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32817\
        );

    \I__6355\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32817\
        );

    \I__6354\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32814\
        );

    \I__6353\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32811\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__32817\,
            I => \N__32808\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__32814\,
            I => \elapsed_time_ns_1_RNIGH4DM1_0_17\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__32811\,
            I => \elapsed_time_ns_1_RNIGH4DM1_0_17\
        );

    \I__6349\ : Odrv4
    port map (
            O => \N__32808\,
            I => \elapsed_time_ns_1_RNIGH4DM1_0_17\
        );

    \I__6348\ : InMux
    port map (
            O => \N__32801\,
            I => \N__32798\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__32798\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9\
        );

    \I__6346\ : CascadeMux
    port map (
            O => \N__32795\,
            I => \N__32791\
        );

    \I__6345\ : InMux
    port map (
            O => \N__32794\,
            I => \N__32788\
        );

    \I__6344\ : InMux
    port map (
            O => \N__32791\,
            I => \N__32785\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__32788\,
            I => \N__32782\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__32785\,
            I => \N__32779\
        );

    \I__6341\ : Odrv4
    port map (
            O => \N__32782\,
            I => \phase_controller_inst1.stoper_tr.N_251\
        );

    \I__6340\ : Odrv4
    port map (
            O => \N__32779\,
            I => \phase_controller_inst1.stoper_tr.N_251\
        );

    \I__6339\ : CascadeMux
    port map (
            O => \N__32774\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\
        );

    \I__6338\ : InMux
    port map (
            O => \N__32771\,
            I => \N__32768\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__32768\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\
        );

    \I__6336\ : InMux
    port map (
            O => \N__32765\,
            I => \N__32760\
        );

    \I__6335\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32755\
        );

    \I__6334\ : InMux
    port map (
            O => \N__32763\,
            I => \N__32755\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__32760\,
            I => \N__32748\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__32755\,
            I => \N__32748\
        );

    \I__6331\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32743\
        );

    \I__6330\ : InMux
    port map (
            O => \N__32753\,
            I => \N__32743\
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__32748\,
            I => \elapsed_time_ns_1_RNI1OL2M1_0_9\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__32743\,
            I => \elapsed_time_ns_1_RNI1OL2M1_0_9\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__32738\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\
        );

    \I__6326\ : CascadeMux
    port map (
            O => \N__32735\,
            I => \N__32731\
        );

    \I__6325\ : InMux
    port map (
            O => \N__32734\,
            I => \N__32727\
        );

    \I__6324\ : InMux
    port map (
            O => \N__32731\,
            I => \N__32724\
        );

    \I__6323\ : InMux
    port map (
            O => \N__32730\,
            I => \N__32721\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__32727\,
            I => \N__32717\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__32724\,
            I => \N__32712\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__32721\,
            I => \N__32712\
        );

    \I__6319\ : InMux
    port map (
            O => \N__32720\,
            I => \N__32709\
        );

    \I__6318\ : Span4Mux_h
    port map (
            O => \N__32717\,
            I => \N__32706\
        );

    \I__6317\ : Odrv4
    port map (
            O => \N__32712\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__32709\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6315\ : Odrv4
    port map (
            O => \N__32706\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6314\ : CascadeMux
    port map (
            O => \N__32699\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\
        );

    \I__6313\ : InMux
    port map (
            O => \N__32696\,
            I => \N__32690\
        );

    \I__6312\ : InMux
    port map (
            O => \N__32695\,
            I => \N__32690\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__32690\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__32687\,
            I => \elapsed_time_ns_1_RNICG2591_0_4_cascade_\
        );

    \I__6309\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32681\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__32681\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2\
        );

    \I__6307\ : CascadeMux
    port map (
            O => \N__32678\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_\
        );

    \I__6306\ : CascadeMux
    port map (
            O => \N__32675\,
            I => \N__32671\
        );

    \I__6305\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32665\
        );

    \I__6304\ : InMux
    port map (
            O => \N__32671\,
            I => \N__32662\
        );

    \I__6303\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32655\
        );

    \I__6302\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32655\
        );

    \I__6301\ : InMux
    port map (
            O => \N__32668\,
            I => \N__32655\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__32665\,
            I => \elapsed_time_ns_1_RNIFG4DM1_0_16\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__32662\,
            I => \elapsed_time_ns_1_RNIFG4DM1_0_16\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__32655\,
            I => \elapsed_time_ns_1_RNIFG4DM1_0_16\
        );

    \I__6297\ : CascadeMux
    port map (
            O => \N__32648\,
            I => \elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_\
        );

    \I__6296\ : InMux
    port map (
            O => \N__32645\,
            I => \N__32642\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__32642\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\
        );

    \I__6294\ : CascadeMux
    port map (
            O => \N__32639\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18_cascade_\
        );

    \I__6293\ : CascadeMux
    port map (
            O => \N__32636\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\
        );

    \I__6292\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32630\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__32630\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\
        );

    \I__6290\ : CascadeMux
    port map (
            O => \N__32627\,
            I => \elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_\
        );

    \I__6289\ : CascadeMux
    port map (
            O => \N__32624\,
            I => \phase_controller_inst1.stoper_tr.N_211_cascade_\
        );

    \I__6288\ : CascadeMux
    port map (
            O => \N__32621\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_\
        );

    \I__6287\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32615\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__32615\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\
        );

    \I__6285\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32605\
        );

    \I__6284\ : InMux
    port map (
            O => \N__32611\,
            I => \N__32605\
        );

    \I__6283\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32602\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__32605\,
            I => \elapsed_time_ns_1_RNIPFL2M1_0_1\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__32602\,
            I => \elapsed_time_ns_1_RNIPFL2M1_0_1\
        );

    \I__6280\ : InMux
    port map (
            O => \N__32597\,
            I => \N__32593\
        );

    \I__6279\ : InMux
    port map (
            O => \N__32596\,
            I => \N__32590\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__32593\,
            I => \N__32587\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__32590\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\
        );

    \I__6276\ : Odrv4
    port map (
            O => \N__32587\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\
        );

    \I__6275\ : CascadeMux
    port map (
            O => \N__32582\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_\
        );

    \I__6274\ : CascadeMux
    port map (
            O => \N__32579\,
            I => \N__32571\
        );

    \I__6273\ : CascadeMux
    port map (
            O => \N__32578\,
            I => \N__32568\
        );

    \I__6272\ : CascadeMux
    port map (
            O => \N__32577\,
            I => \N__32564\
        );

    \I__6271\ : CascadeMux
    port map (
            O => \N__32576\,
            I => \N__32561\
        );

    \I__6270\ : CascadeMux
    port map (
            O => \N__32575\,
            I => \N__32555\
        );

    \I__6269\ : CascadeMux
    port map (
            O => \N__32574\,
            I => \N__32552\
        );

    \I__6268\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32548\
        );

    \I__6267\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32545\
        );

    \I__6266\ : InMux
    port map (
            O => \N__32567\,
            I => \N__32542\
        );

    \I__6265\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32539\
        );

    \I__6264\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32534\
        );

    \I__6263\ : InMux
    port map (
            O => \N__32560\,
            I => \N__32534\
        );

    \I__6262\ : InMux
    port map (
            O => \N__32559\,
            I => \N__32523\
        );

    \I__6261\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32523\
        );

    \I__6260\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32523\
        );

    \I__6259\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32523\
        );

    \I__6258\ : InMux
    port map (
            O => \N__32551\,
            I => \N__32523\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__32548\,
            I => \N__32518\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__32545\,
            I => \N__32518\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__32542\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__32539\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__32534\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__32523\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__6251\ : Odrv12
    port map (
            O => \N__32518\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__6250\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32498\
        );

    \I__6249\ : InMux
    port map (
            O => \N__32506\,
            I => \N__32498\
        );

    \I__6248\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32498\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__32498\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2\
        );

    \I__6246\ : CascadeMux
    port map (
            O => \N__32495\,
            I => \N__32491\
        );

    \I__6245\ : InMux
    port map (
            O => \N__32494\,
            I => \N__32488\
        );

    \I__6244\ : InMux
    port map (
            O => \N__32491\,
            I => \N__32485\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__32488\,
            I => \N__32479\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__32485\,
            I => \N__32479\
        );

    \I__6241\ : InMux
    port map (
            O => \N__32484\,
            I => \N__32476\
        );

    \I__6240\ : Odrv4
    port map (
            O => \N__32479\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__32476\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__6238\ : CEMux
    port map (
            O => \N__32471\,
            I => \N__32466\
        );

    \I__6237\ : CEMux
    port map (
            O => \N__32470\,
            I => \N__32463\
        );

    \I__6236\ : CEMux
    port map (
            O => \N__32469\,
            I => \N__32459\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__32466\,
            I => \N__32454\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__32463\,
            I => \N__32454\
        );

    \I__6233\ : CEMux
    port map (
            O => \N__32462\,
            I => \N__32451\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__32459\,
            I => \N__32448\
        );

    \I__6231\ : Span4Mux_v
    port map (
            O => \N__32454\,
            I => \N__32445\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__32451\,
            I => \N__32442\
        );

    \I__6229\ : Span4Mux_v
    port map (
            O => \N__32448\,
            I => \N__32435\
        );

    \I__6228\ : Span4Mux_h
    port map (
            O => \N__32445\,
            I => \N__32435\
        );

    \I__6227\ : Span4Mux_h
    port map (
            O => \N__32442\,
            I => \N__32435\
        );

    \I__6226\ : Span4Mux_h
    port map (
            O => \N__32435\,
            I => \N__32432\
        );

    \I__6225\ : Odrv4
    port map (
            O => \N__32432\,
            I => \delay_measurement_inst.delay_hc_timer.N_433_i\
        );

    \I__6224\ : InMux
    port map (
            O => \N__32429\,
            I => \N__32425\
        );

    \I__6223\ : InMux
    port map (
            O => \N__32428\,
            I => \N__32420\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__32425\,
            I => \N__32417\
        );

    \I__6221\ : InMux
    port map (
            O => \N__32424\,
            I => \N__32412\
        );

    \I__6220\ : InMux
    port map (
            O => \N__32423\,
            I => \N__32412\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__32420\,
            I => \N__32407\
        );

    \I__6218\ : Span12Mux_s7_v
    port map (
            O => \N__32417\,
            I => \N__32407\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__32412\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6216\ : Odrv12
    port map (
            O => \N__32407\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6215\ : IoInMux
    port map (
            O => \N__32402\,
            I => \N__32399\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__32399\,
            I => \N__32396\
        );

    \I__6213\ : Odrv12
    port map (
            O => \N__32396\,
            I => \current_shift_inst.timer_s1.N_166_i\
        );

    \I__6212\ : CascadeMux
    port map (
            O => \N__32393\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_\
        );

    \I__6211\ : CascadeMux
    port map (
            O => \N__32390\,
            I => \elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_\
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__32387\,
            I => \N__32383\
        );

    \I__6209\ : CascadeMux
    port map (
            O => \N__32386\,
            I => \N__32379\
        );

    \I__6208\ : InMux
    port map (
            O => \N__32383\,
            I => \N__32376\
        );

    \I__6207\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32373\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32379\,
            I => \N__32370\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__32376\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__32373\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__32370\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6\
        );

    \I__6202\ : InMux
    port map (
            O => \N__32363\,
            I => \N__32359\
        );

    \I__6201\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32356\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__32359\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__32356\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__32351\,
            I => \N__32348\
        );

    \I__6197\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32343\
        );

    \I__6196\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32340\
        );

    \I__6195\ : InMux
    port map (
            O => \N__32346\,
            I => \N__32337\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__32343\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__32340\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__32337\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__6191\ : InMux
    port map (
            O => \N__32330\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__6190\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32322\
        );

    \I__6189\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32317\
        );

    \I__6188\ : InMux
    port map (
            O => \N__32325\,
            I => \N__32317\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__32322\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__32317\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__6185\ : InMux
    port map (
            O => \N__32312\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__6184\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32304\
        );

    \I__6183\ : InMux
    port map (
            O => \N__32308\,
            I => \N__32299\
        );

    \I__6182\ : InMux
    port map (
            O => \N__32307\,
            I => \N__32299\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__32304\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__32299\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__6179\ : InMux
    port map (
            O => \N__32294\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__6178\ : CascadeMux
    port map (
            O => \N__32291\,
            I => \N__32287\
        );

    \I__6177\ : CascadeMux
    port map (
            O => \N__32290\,
            I => \N__32284\
        );

    \I__6176\ : InMux
    port map (
            O => \N__32287\,
            I => \N__32280\
        );

    \I__6175\ : InMux
    port map (
            O => \N__32284\,
            I => \N__32277\
        );

    \I__6174\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32274\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__32280\,
            I => \N__32271\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__32277\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__32274\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__32271\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__6169\ : InMux
    port map (
            O => \N__32264\,
            I => \bfn_13_24_0_\
        );

    \I__6168\ : CascadeMux
    port map (
            O => \N__32261\,
            I => \N__32257\
        );

    \I__6167\ : CascadeMux
    port map (
            O => \N__32260\,
            I => \N__32254\
        );

    \I__6166\ : InMux
    port map (
            O => \N__32257\,
            I => \N__32250\
        );

    \I__6165\ : InMux
    port map (
            O => \N__32254\,
            I => \N__32247\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32253\,
            I => \N__32244\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__32250\,
            I => \N__32241\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__32247\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__32244\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__6160\ : Odrv4
    port map (
            O => \N__32241\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__6159\ : InMux
    port map (
            O => \N__32234\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__6158\ : CascadeMux
    port map (
            O => \N__32231\,
            I => \N__32228\
        );

    \I__6157\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32223\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32227\,
            I => \N__32220\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32226\,
            I => \N__32217\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__32223\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__32220\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__32217\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__6151\ : InMux
    port map (
            O => \N__32210\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__6150\ : CascadeMux
    port map (
            O => \N__32207\,
            I => \N__32204\
        );

    \I__6149\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32199\
        );

    \I__6148\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32196\
        );

    \I__6147\ : InMux
    port map (
            O => \N__32202\,
            I => \N__32193\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__32199\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__32196\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__32193\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__6143\ : InMux
    port map (
            O => \N__32186\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32183\,
            I => \N__32179\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32176\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__32179\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__32176\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__6138\ : InMux
    port map (
            O => \N__32171\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__6137\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32130\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32130\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32130\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32130\
        );

    \I__6133\ : InMux
    port map (
            O => \N__32164\,
            I => \N__32125\
        );

    \I__6132\ : InMux
    port map (
            O => \N__32163\,
            I => \N__32125\
        );

    \I__6131\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32116\
        );

    \I__6130\ : InMux
    port map (
            O => \N__32161\,
            I => \N__32116\
        );

    \I__6129\ : InMux
    port map (
            O => \N__32160\,
            I => \N__32116\
        );

    \I__6128\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32116\
        );

    \I__6127\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32107\
        );

    \I__6126\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32107\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32107\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32155\,
            I => \N__32107\
        );

    \I__6123\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32098\
        );

    \I__6122\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32098\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32152\,
            I => \N__32098\
        );

    \I__6120\ : InMux
    port map (
            O => \N__32151\,
            I => \N__32098\
        );

    \I__6119\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32089\
        );

    \I__6118\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32089\
        );

    \I__6117\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32089\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32089\
        );

    \I__6115\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32080\
        );

    \I__6114\ : InMux
    port map (
            O => \N__32145\,
            I => \N__32080\
        );

    \I__6113\ : InMux
    port map (
            O => \N__32144\,
            I => \N__32080\
        );

    \I__6112\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32080\
        );

    \I__6111\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32071\
        );

    \I__6110\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32071\
        );

    \I__6109\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32071\
        );

    \I__6108\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32071\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__32130\,
            I => \N__32068\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__32125\,
            I => \N__32057\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__32116\,
            I => \N__32057\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__32107\,
            I => \N__32057\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__32098\,
            I => \N__32057\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__32089\,
            I => \N__32057\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__32080\,
            I => \N__32052\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__32071\,
            I => \N__32052\
        );

    \I__6099\ : Span4Mux_v
    port map (
            O => \N__32068\,
            I => \N__32047\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__32057\,
            I => \N__32047\
        );

    \I__6097\ : Span4Mux_h
    port map (
            O => \N__32052\,
            I => \N__32044\
        );

    \I__6096\ : Odrv4
    port map (
            O => \N__32047\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__32044\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__6094\ : InMux
    port map (
            O => \N__32039\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__6093\ : InMux
    port map (
            O => \N__32036\,
            I => \N__32032\
        );

    \I__6092\ : InMux
    port map (
            O => \N__32035\,
            I => \N__32029\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__32032\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__32029\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__6089\ : CascadeMux
    port map (
            O => \N__32024\,
            I => \N__32021\
        );

    \I__6088\ : InMux
    port map (
            O => \N__32021\,
            I => \N__32016\
        );

    \I__6087\ : InMux
    port map (
            O => \N__32020\,
            I => \N__32013\
        );

    \I__6086\ : InMux
    port map (
            O => \N__32019\,
            I => \N__32010\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__32016\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32013\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__32010\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__6082\ : InMux
    port map (
            O => \N__32003\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__6081\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31995\
        );

    \I__6080\ : InMux
    port map (
            O => \N__31999\,
            I => \N__31990\
        );

    \I__6079\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31990\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__31995\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__31990\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__6076\ : InMux
    port map (
            O => \N__31985\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__6075\ : InMux
    port map (
            O => \N__31982\,
            I => \N__31977\
        );

    \I__6074\ : InMux
    port map (
            O => \N__31981\,
            I => \N__31972\
        );

    \I__6073\ : InMux
    port map (
            O => \N__31980\,
            I => \N__31972\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__31977\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__31972\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__6070\ : InMux
    port map (
            O => \N__31967\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__6069\ : CascadeMux
    port map (
            O => \N__31964\,
            I => \N__31961\
        );

    \I__6068\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31957\
        );

    \I__6067\ : CascadeMux
    port map (
            O => \N__31960\,
            I => \N__31954\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__31957\,
            I => \N__31950\
        );

    \I__6065\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31947\
        );

    \I__6064\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31944\
        );

    \I__6063\ : Span4Mux_h
    port map (
            O => \N__31950\,
            I => \N__31941\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__31947\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__31944\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__31941\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__6059\ : InMux
    port map (
            O => \N__31934\,
            I => \bfn_13_23_0_\
        );

    \I__6058\ : CascadeMux
    port map (
            O => \N__31931\,
            I => \N__31927\
        );

    \I__6057\ : CascadeMux
    port map (
            O => \N__31930\,
            I => \N__31924\
        );

    \I__6056\ : InMux
    port map (
            O => \N__31927\,
            I => \N__31920\
        );

    \I__6055\ : InMux
    port map (
            O => \N__31924\,
            I => \N__31917\
        );

    \I__6054\ : InMux
    port map (
            O => \N__31923\,
            I => \N__31914\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__31920\,
            I => \N__31911\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__31917\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__31914\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__6050\ : Odrv4
    port map (
            O => \N__31911\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__6049\ : InMux
    port map (
            O => \N__31904\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__6048\ : InMux
    port map (
            O => \N__31901\,
            I => \N__31897\
        );

    \I__6047\ : CascadeMux
    port map (
            O => \N__31900\,
            I => \N__31894\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__31897\,
            I => \N__31890\
        );

    \I__6045\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31887\
        );

    \I__6044\ : InMux
    port map (
            O => \N__31893\,
            I => \N__31884\
        );

    \I__6043\ : Span4Mux_h
    port map (
            O => \N__31890\,
            I => \N__31881\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__31887\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__31884\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__31881\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__6039\ : InMux
    port map (
            O => \N__31874\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__6038\ : CascadeMux
    port map (
            O => \N__31871\,
            I => \N__31868\
        );

    \I__6037\ : InMux
    port map (
            O => \N__31868\,
            I => \N__31863\
        );

    \I__6036\ : InMux
    port map (
            O => \N__31867\,
            I => \N__31860\
        );

    \I__6035\ : InMux
    port map (
            O => \N__31866\,
            I => \N__31857\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__31863\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__31860\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__31857\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__6031\ : InMux
    port map (
            O => \N__31850\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__31847\,
            I => \N__31844\
        );

    \I__6029\ : InMux
    port map (
            O => \N__31844\,
            I => \N__31839\
        );

    \I__6028\ : InMux
    port map (
            O => \N__31843\,
            I => \N__31836\
        );

    \I__6027\ : InMux
    port map (
            O => \N__31842\,
            I => \N__31833\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__31839\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__31836\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__31833\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__6023\ : InMux
    port map (
            O => \N__31826\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__6022\ : InMux
    port map (
            O => \N__31823\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__6021\ : CascadeMux
    port map (
            O => \N__31820\,
            I => \N__31817\
        );

    \I__6020\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31812\
        );

    \I__6019\ : InMux
    port map (
            O => \N__31816\,
            I => \N__31809\
        );

    \I__6018\ : InMux
    port map (
            O => \N__31815\,
            I => \N__31806\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__31812\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__31809\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__31806\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__6014\ : InMux
    port map (
            O => \N__31799\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__6013\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31791\
        );

    \I__6012\ : InMux
    port map (
            O => \N__31795\,
            I => \N__31786\
        );

    \I__6011\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31786\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__31791\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__31786\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__6008\ : InMux
    port map (
            O => \N__31781\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__6007\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31773\
        );

    \I__6006\ : InMux
    port map (
            O => \N__31777\,
            I => \N__31768\
        );

    \I__6005\ : InMux
    port map (
            O => \N__31776\,
            I => \N__31768\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__31773\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__31768\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__6002\ : InMux
    port map (
            O => \N__31763\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__31760\,
            I => \N__31756\
        );

    \I__6000\ : CascadeMux
    port map (
            O => \N__31759\,
            I => \N__31753\
        );

    \I__5999\ : InMux
    port map (
            O => \N__31756\,
            I => \N__31749\
        );

    \I__5998\ : InMux
    port map (
            O => \N__31753\,
            I => \N__31746\
        );

    \I__5997\ : InMux
    port map (
            O => \N__31752\,
            I => \N__31743\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__31749\,
            I => \N__31740\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__31746\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__31743\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__5993\ : Odrv4
    port map (
            O => \N__31740\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__5992\ : InMux
    port map (
            O => \N__31733\,
            I => \bfn_13_22_0_\
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__31730\,
            I => \N__31726\
        );

    \I__5990\ : CascadeMux
    port map (
            O => \N__31729\,
            I => \N__31723\
        );

    \I__5989\ : InMux
    port map (
            O => \N__31726\,
            I => \N__31719\
        );

    \I__5988\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31716\
        );

    \I__5987\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31713\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__31719\,
            I => \N__31710\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__31716\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__31713\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__5983\ : Odrv4
    port map (
            O => \N__31710\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__5982\ : InMux
    port map (
            O => \N__31703\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__31700\,
            I => \N__31697\
        );

    \I__5980\ : InMux
    port map (
            O => \N__31697\,
            I => \N__31692\
        );

    \I__5979\ : InMux
    port map (
            O => \N__31696\,
            I => \N__31689\
        );

    \I__5978\ : InMux
    port map (
            O => \N__31695\,
            I => \N__31686\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__31692\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__31689\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__31686\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__5974\ : InMux
    port map (
            O => \N__31679\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__5973\ : CascadeMux
    port map (
            O => \N__31676\,
            I => \N__31673\
        );

    \I__5972\ : InMux
    port map (
            O => \N__31673\,
            I => \N__31668\
        );

    \I__5971\ : InMux
    port map (
            O => \N__31672\,
            I => \N__31665\
        );

    \I__5970\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31662\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__31668\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__31665\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__31662\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__5966\ : InMux
    port map (
            O => \N__31655\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__5965\ : CascadeMux
    port map (
            O => \N__31652\,
            I => \N__31649\
        );

    \I__5964\ : InMux
    port map (
            O => \N__31649\,
            I => \N__31644\
        );

    \I__5963\ : InMux
    port map (
            O => \N__31648\,
            I => \N__31641\
        );

    \I__5962\ : InMux
    port map (
            O => \N__31647\,
            I => \N__31638\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__31644\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__31641\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__31638\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__5958\ : InMux
    port map (
            O => \N__31631\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__5957\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31625\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__31625\,
            I => \N__31622\
        );

    \I__5955\ : Span4Mux_h
    port map (
            O => \N__31622\,
            I => \N__31619\
        );

    \I__5954\ : Span4Mux_h
    port map (
            O => \N__31619\,
            I => \N__31616\
        );

    \I__5953\ : Odrv4
    port map (
            O => \N__31616\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__5952\ : InMux
    port map (
            O => \N__31613\,
            I => \bfn_13_21_0_\
        );

    \I__5951\ : InMux
    port map (
            O => \N__31610\,
            I => \N__31607\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__31607\,
            I => \N__31604\
        );

    \I__5949\ : Span4Mux_h
    port map (
            O => \N__31604\,
            I => \N__31600\
        );

    \I__5948\ : CascadeMux
    port map (
            O => \N__31603\,
            I => \N__31597\
        );

    \I__5947\ : Span4Mux_h
    port map (
            O => \N__31600\,
            I => \N__31593\
        );

    \I__5946\ : InMux
    port map (
            O => \N__31597\,
            I => \N__31590\
        );

    \I__5945\ : InMux
    port map (
            O => \N__31596\,
            I => \N__31587\
        );

    \I__5944\ : Odrv4
    port map (
            O => \N__31593\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__31590\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__31587\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__5941\ : InMux
    port map (
            O => \N__31580\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__5940\ : CascadeMux
    port map (
            O => \N__31577\,
            I => \N__31574\
        );

    \I__5939\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31569\
        );

    \I__5938\ : InMux
    port map (
            O => \N__31573\,
            I => \N__31566\
        );

    \I__5937\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31563\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__31569\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__31566\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__31563\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__5933\ : InMux
    port map (
            O => \N__31556\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__5932\ : CascadeMux
    port map (
            O => \N__31553\,
            I => \N__31550\
        );

    \I__5931\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31545\
        );

    \I__5930\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31542\
        );

    \I__5929\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31539\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__31545\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__31542\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__31539\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__5925\ : InMux
    port map (
            O => \N__31532\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__5924\ : CascadeMux
    port map (
            O => \N__31529\,
            I => \N__31526\
        );

    \I__5923\ : InMux
    port map (
            O => \N__31526\,
            I => \N__31521\
        );

    \I__5922\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31518\
        );

    \I__5921\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31515\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__31521\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__31518\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__31515\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__5917\ : InMux
    port map (
            O => \N__31508\,
            I => \N__31504\
        );

    \I__5916\ : CascadeMux
    port map (
            O => \N__31507\,
            I => \N__31499\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__31504\,
            I => \N__31496\
        );

    \I__5914\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31489\
        );

    \I__5913\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31489\
        );

    \I__5912\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31489\
        );

    \I__5911\ : Span4Mux_v
    port map (
            O => \N__31496\,
            I => \N__31486\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__31489\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__5909\ : Odrv4
    port map (
            O => \N__31486\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__31481\,
            I => \N__31477\
        );

    \I__5907\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31466\
        );

    \I__5906\ : InMux
    port map (
            O => \N__31477\,
            I => \N__31466\
        );

    \I__5905\ : InMux
    port map (
            O => \N__31476\,
            I => \N__31466\
        );

    \I__5904\ : InMux
    port map (
            O => \N__31475\,
            I => \N__31466\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__31466\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__5902\ : CascadeMux
    port map (
            O => \N__31463\,
            I => \N__31460\
        );

    \I__5901\ : InMux
    port map (
            O => \N__31460\,
            I => \N__31456\
        );

    \I__5900\ : InMux
    port map (
            O => \N__31459\,
            I => \N__31452\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__31456\,
            I => \N__31449\
        );

    \I__5898\ : InMux
    port map (
            O => \N__31455\,
            I => \N__31445\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__31452\,
            I => \N__31442\
        );

    \I__5896\ : Span4Mux_h
    port map (
            O => \N__31449\,
            I => \N__31439\
        );

    \I__5895\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31436\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__31445\,
            I => \N__31431\
        );

    \I__5893\ : Span4Mux_h
    port map (
            O => \N__31442\,
            I => \N__31431\
        );

    \I__5892\ : Span4Mux_h
    port map (
            O => \N__31439\,
            I => \N__31428\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__31436\,
            I => \N__31423\
        );

    \I__5890\ : Span4Mux_v
    port map (
            O => \N__31431\,
            I => \N__31423\
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__31428\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__31423\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5887\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31415\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__31415\,
            I => \N__31412\
        );

    \I__5885\ : Odrv12
    port map (
            O => \N__31412\,
            I => \current_shift_inst.PI_CTRL.integrator_i_30\
        );

    \I__5884\ : InMux
    port map (
            O => \N__31409\,
            I => \N__31405\
        );

    \I__5883\ : InMux
    port map (
            O => \N__31408\,
            I => \N__31402\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__31405\,
            I => \N__31398\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__31402\,
            I => \N__31395\
        );

    \I__5880\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31392\
        );

    \I__5879\ : Span4Mux_v
    port map (
            O => \N__31398\,
            I => \N__31387\
        );

    \I__5878\ : Span4Mux_v
    port map (
            O => \N__31395\,
            I => \N__31384\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__31392\,
            I => \N__31381\
        );

    \I__5876\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31376\
        );

    \I__5875\ : InMux
    port map (
            O => \N__31390\,
            I => \N__31376\
        );

    \I__5874\ : Span4Mux_v
    port map (
            O => \N__31387\,
            I => \N__31369\
        );

    \I__5873\ : Span4Mux_h
    port map (
            O => \N__31384\,
            I => \N__31369\
        );

    \I__5872\ : Span4Mux_v
    port map (
            O => \N__31381\,
            I => \N__31369\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__31376\,
            I => \N__31366\
        );

    \I__5870\ : Odrv4
    port map (
            O => \N__31369\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5869\ : Odrv12
    port map (
            O => \N__31366\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5868\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31358\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__31358\,
            I => \N__31355\
        );

    \I__5866\ : Odrv12
    port map (
            O => \N__31355\,
            I => \current_shift_inst.PI_CTRL.integrator_i_27\
        );

    \I__5865\ : CascadeMux
    port map (
            O => \N__31352\,
            I => \N__31349\
        );

    \I__5864\ : InMux
    port map (
            O => \N__31349\,
            I => \N__31346\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__31346\,
            I => \N__31342\
        );

    \I__5862\ : CascadeMux
    port map (
            O => \N__31345\,
            I => \N__31339\
        );

    \I__5861\ : Span4Mux_v
    port map (
            O => \N__31342\,
            I => \N__31335\
        );

    \I__5860\ : InMux
    port map (
            O => \N__31339\,
            I => \N__31329\
        );

    \I__5859\ : InMux
    port map (
            O => \N__31338\,
            I => \N__31329\
        );

    \I__5858\ : Span4Mux_h
    port map (
            O => \N__31335\,
            I => \N__31326\
        );

    \I__5857\ : InMux
    port map (
            O => \N__31334\,
            I => \N__31323\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__31329\,
            I => \N__31320\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__31326\,
            I => \N__31315\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__31323\,
            I => \N__31315\
        );

    \I__5853\ : Span4Mux_h
    port map (
            O => \N__31320\,
            I => \N__31312\
        );

    \I__5852\ : Odrv4
    port map (
            O => \N__31315\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__5851\ : Odrv4
    port map (
            O => \N__31312\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__5850\ : InMux
    port map (
            O => \N__31307\,
            I => \N__31304\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__31304\,
            I => \N__31301\
        );

    \I__5848\ : Odrv12
    port map (
            O => \N__31301\,
            I => \current_shift_inst.PI_CTRL.integrator_i_28\
        );

    \I__5847\ : CascadeMux
    port map (
            O => \N__31298\,
            I => \N__31295\
        );

    \I__5846\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31291\
        );

    \I__5845\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31288\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__31291\,
            I => \N__31282\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__31288\,
            I => \N__31282\
        );

    \I__5842\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31279\
        );

    \I__5841\ : Span4Mux_h
    port map (
            O => \N__31282\,
            I => \N__31276\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__31279\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__5839\ : Odrv4
    port map (
            O => \N__31276\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__5838\ : InMux
    port map (
            O => \N__31271\,
            I => \N__31262\
        );

    \I__5837\ : InMux
    port map (
            O => \N__31270\,
            I => \N__31262\
        );

    \I__5836\ : InMux
    port map (
            O => \N__31269\,
            I => \N__31262\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__31262\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__5834\ : CascadeMux
    port map (
            O => \N__31259\,
            I => \phase_controller_inst2.time_passed_RNI9M3O_cascade_\
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__31256\,
            I => \N__31249\
        );

    \I__5832\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31242\
        );

    \I__5831\ : InMux
    port map (
            O => \N__31254\,
            I => \N__31242\
        );

    \I__5830\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31242\
        );

    \I__5829\ : CascadeMux
    port map (
            O => \N__31252\,
            I => \N__31239\
        );

    \I__5828\ : InMux
    port map (
            O => \N__31249\,
            I => \N__31235\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__31242\,
            I => \N__31232\
        );

    \I__5826\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31229\
        );

    \I__5825\ : InMux
    port map (
            O => \N__31238\,
            I => \N__31226\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__31235\,
            I => \N__31221\
        );

    \I__5823\ : Span4Mux_v
    port map (
            O => \N__31232\,
            I => \N__31221\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__31229\,
            I => \N__31216\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__31226\,
            I => \N__31216\
        );

    \I__5820\ : Odrv4
    port map (
            O => \N__31221\,
            I => state_3
        );

    \I__5819\ : Odrv4
    port map (
            O => \N__31216\,
            I => state_3
        );

    \I__5818\ : IoInMux
    port map (
            O => \N__31211\,
            I => \N__31208\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__31208\,
            I => \N__31205\
        );

    \I__5816\ : Span4Mux_s3_v
    port map (
            O => \N__31205\,
            I => \N__31202\
        );

    \I__5815\ : Sp12to4
    port map (
            O => \N__31202\,
            I => \N__31199\
        );

    \I__5814\ : Span12Mux_h
    port map (
            O => \N__31199\,
            I => \N__31196\
        );

    \I__5813\ : Span12Mux_v
    port map (
            O => \N__31196\,
            I => \N__31191\
        );

    \I__5812\ : InMux
    port map (
            O => \N__31195\,
            I => \N__31186\
        );

    \I__5811\ : InMux
    port map (
            O => \N__31194\,
            I => \N__31186\
        );

    \I__5810\ : Odrv12
    port map (
            O => \N__31191\,
            I => s1_phy_c
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__31186\,
            I => s1_phy_c
        );

    \I__5808\ : InMux
    port map (
            O => \N__31181\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__5807\ : InMux
    port map (
            O => \N__31178\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__5806\ : InMux
    port map (
            O => \N__31175\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__5805\ : InMux
    port map (
            O => \N__31172\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31169\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__5803\ : InMux
    port map (
            O => \N__31166\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__5802\ : InMux
    port map (
            O => \N__31163\,
            I => \bfn_13_13_0_\
        );

    \I__5801\ : InMux
    port map (
            O => \N__31160\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__5800\ : InMux
    port map (
            O => \N__31157\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__5799\ : InMux
    port map (
            O => \N__31154\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__5798\ : InMux
    port map (
            O => \N__31151\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__5797\ : InMux
    port map (
            O => \N__31148\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__5796\ : InMux
    port map (
            O => \N__31145\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__5795\ : InMux
    port map (
            O => \N__31142\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__5794\ : InMux
    port map (
            O => \N__31139\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__5793\ : InMux
    port map (
            O => \N__31136\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__5792\ : InMux
    port map (
            O => \N__31133\,
            I => \bfn_13_12_0_\
        );

    \I__5791\ : InMux
    port map (
            O => \N__31130\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__5790\ : CascadeMux
    port map (
            O => \N__31127\,
            I => \N__31123\
        );

    \I__5789\ : InMux
    port map (
            O => \N__31126\,
            I => \N__31120\
        );

    \I__5788\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31117\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__31120\,
            I => \N__31114\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__31117\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__31114\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\
        );

    \I__5784\ : CascadeMux
    port map (
            O => \N__31109\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_\
        );

    \I__5783\ : CascadeMux
    port map (
            O => \N__31106\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_\
        );

    \I__5782\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31094\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31094\
        );

    \I__5780\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31094\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__31094\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2\
        );

    \I__5778\ : CascadeMux
    port map (
            O => \N__31091\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_\
        );

    \I__5777\ : CascadeMux
    port map (
            O => \N__31088\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_\
        );

    \I__5776\ : CascadeMux
    port map (
            O => \N__31085\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19_cascade_\
        );

    \I__5775\ : CascadeMux
    port map (
            O => \N__31082\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_\
        );

    \I__5774\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31075\
        );

    \I__5773\ : InMux
    port map (
            O => \N__31078\,
            I => \N__31070\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__31075\,
            I => \N__31067\
        );

    \I__5771\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31064\
        );

    \I__5770\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31061\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__31070\,
            I => \N__31056\
        );

    \I__5768\ : Span12Mux_s9_v
    port map (
            O => \N__31067\,
            I => \N__31056\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__31064\,
            I => \N__31053\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__31061\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__5765\ : Odrv12
    port map (
            O => \N__31056\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__31053\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__5763\ : IoInMux
    port map (
            O => \N__31046\,
            I => \N__31043\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__31043\,
            I => \N__31040\
        );

    \I__5761\ : Span4Mux_s1_v
    port map (
            O => \N__31040\,
            I => \N__31037\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__31037\,
            I => s2_phy_c
        );

    \I__5759\ : IoInMux
    port map (
            O => \N__31034\,
            I => \N__31031\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__31031\,
            I => \N__31028\
        );

    \I__5757\ : Span4Mux_s0_v
    port map (
            O => \N__31028\,
            I => \N__31025\
        );

    \I__5756\ : Odrv4
    port map (
            O => \N__31025\,
            I => \pll_inst.red_c_i\
        );

    \I__5755\ : InMux
    port map (
            O => \N__31022\,
            I => \N__31019\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__31019\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1\
        );

    \I__5753\ : InMux
    port map (
            O => \N__31016\,
            I => \N__31012\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__31015\,
            I => \N__31009\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__31012\,
            I => \N__31006\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31009\,
            I => \N__31003\
        );

    \I__5749\ : Odrv4
    port map (
            O => \N__31006\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__31003\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__5747\ : InMux
    port map (
            O => \N__30998\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__30995\,
            I => \N__30992\
        );

    \I__5745\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30989\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__30989\,
            I => \N__30986\
        );

    \I__5743\ : Span4Mux_v
    port map (
            O => \N__30986\,
            I => \N__30982\
        );

    \I__5742\ : InMux
    port map (
            O => \N__30985\,
            I => \N__30979\
        );

    \I__5741\ : Odrv4
    port map (
            O => \N__30982\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__30979\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__5739\ : InMux
    port map (
            O => \N__30974\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__30971\,
            I => \N__30968\
        );

    \I__5737\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30965\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__30965\,
            I => \N__30962\
        );

    \I__5735\ : Span4Mux_v
    port map (
            O => \N__30962\,
            I => \N__30958\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30961\,
            I => \N__30955\
        );

    \I__5733\ : Odrv4
    port map (
            O => \N__30958\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__30955\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5731\ : InMux
    port map (
            O => \N__30950\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__5730\ : InMux
    port map (
            O => \N__30947\,
            I => \N__30944\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__30944\,
            I => \N__30941\
        );

    \I__5728\ : Span4Mux_h
    port map (
            O => \N__30941\,
            I => \N__30937\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30940\,
            I => \N__30934\
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__30937\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__30934\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__5724\ : InMux
    port map (
            O => \N__30929\,
            I => \bfn_12_23_0_\
        );

    \I__5723\ : InMux
    port map (
            O => \N__30926\,
            I => \N__30923\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__30923\,
            I => \N__30920\
        );

    \I__5721\ : Span4Mux_h
    port map (
            O => \N__30920\,
            I => \N__30916\
        );

    \I__5720\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30913\
        );

    \I__5719\ : Odrv4
    port map (
            O => \N__30916\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__30913\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__5717\ : InMux
    port map (
            O => \N__30908\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__5716\ : CascadeMux
    port map (
            O => \N__30905\,
            I => \N__30902\
        );

    \I__5715\ : InMux
    port map (
            O => \N__30902\,
            I => \N__30899\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__30899\,
            I => \N__30896\
        );

    \I__5713\ : Span4Mux_v
    port map (
            O => \N__30896\,
            I => \N__30892\
        );

    \I__5712\ : InMux
    port map (
            O => \N__30895\,
            I => \N__30889\
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__30892\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__30889\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__5709\ : InMux
    port map (
            O => \N__30884\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__5708\ : InMux
    port map (
            O => \N__30881\,
            I => \N__30878\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__30878\,
            I => \N__30875\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__30875\,
            I => \N__30871\
        );

    \I__5705\ : InMux
    port map (
            O => \N__30874\,
            I => \N__30868\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__30871\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__30868\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__5702\ : InMux
    port map (
            O => \N__30863\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__5701\ : InMux
    port map (
            O => \N__30860\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__5700\ : CascadeMux
    port map (
            O => \N__30857\,
            I => \N__30851\
        );

    \I__5699\ : InMux
    port map (
            O => \N__30856\,
            I => \N__30845\
        );

    \I__5698\ : InMux
    port map (
            O => \N__30855\,
            I => \N__30845\
        );

    \I__5697\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30842\
        );

    \I__5696\ : InMux
    port map (
            O => \N__30851\,
            I => \N__30838\
        );

    \I__5695\ : InMux
    port map (
            O => \N__30850\,
            I => \N__30835\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__30845\,
            I => \N__30830\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__30842\,
            I => \N__30830\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30841\,
            I => \N__30827\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30824\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__30835\,
            I => \N__30821\
        );

    \I__5689\ : Span4Mux_h
    port map (
            O => \N__30830\,
            I => \N__30816\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__30827\,
            I => \N__30816\
        );

    \I__5687\ : Span4Mux_v
    port map (
            O => \N__30824\,
            I => \N__30813\
        );

    \I__5686\ : Span4Mux_v
    port map (
            O => \N__30821\,
            I => \N__30810\
        );

    \I__5685\ : Span4Mux_v
    port map (
            O => \N__30816\,
            I => \N__30807\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__30813\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__5683\ : Odrv4
    port map (
            O => \N__30810\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__5682\ : Odrv4
    port map (
            O => \N__30807\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__5681\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30796\
        );

    \I__5680\ : CascadeMux
    port map (
            O => \N__30799\,
            I => \N__30792\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__30796\,
            I => \N__30787\
        );

    \I__5678\ : InMux
    port map (
            O => \N__30795\,
            I => \N__30782\
        );

    \I__5677\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30782\
        );

    \I__5676\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30777\
        );

    \I__5675\ : InMux
    port map (
            O => \N__30790\,
            I => \N__30777\
        );

    \I__5674\ : Span4Mux_v
    port map (
            O => \N__30787\,
            I => \N__30774\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__30782\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__30777\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5671\ : Odrv4
    port map (
            O => \N__30774\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__30767\,
            I => \N__30764\
        );

    \I__5669\ : InMux
    port map (
            O => \N__30764\,
            I => \N__30760\
        );

    \I__5668\ : CascadeMux
    port map (
            O => \N__30763\,
            I => \N__30757\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__30760\,
            I => \N__30754\
        );

    \I__5666\ : InMux
    port map (
            O => \N__30757\,
            I => \N__30751\
        );

    \I__5665\ : Span4Mux_h
    port map (
            O => \N__30754\,
            I => \N__30747\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__30751\,
            I => \N__30744\
        );

    \I__5663\ : InMux
    port map (
            O => \N__30750\,
            I => \N__30741\
        );

    \I__5662\ : Odrv4
    port map (
            O => \N__30747\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__30744\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__30741\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__5659\ : InMux
    port map (
            O => \N__30734\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__5658\ : InMux
    port map (
            O => \N__30731\,
            I => \N__30728\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__30728\,
            I => \N__30724\
        );

    \I__5656\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30721\
        );

    \I__5655\ : Span4Mux_h
    port map (
            O => \N__30724\,
            I => \N__30717\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__30721\,
            I => \N__30714\
        );

    \I__5653\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30711\
        );

    \I__5652\ : Odrv4
    port map (
            O => \N__30717\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__30714\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__30711\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__5649\ : InMux
    port map (
            O => \N__30704\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__30701\,
            I => \N__30698\
        );

    \I__5647\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30695\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__30695\,
            I => \N__30692\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__30692\,
            I => \N__30688\
        );

    \I__5644\ : InMux
    port map (
            O => \N__30691\,
            I => \N__30685\
        );

    \I__5643\ : Span4Mux_h
    port map (
            O => \N__30688\,
            I => \N__30681\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__30685\,
            I => \N__30678\
        );

    \I__5641\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30675\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__30681\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__5639\ : Odrv4
    port map (
            O => \N__30678\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__30675\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__5637\ : InMux
    port map (
            O => \N__30668\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__5636\ : CascadeMux
    port map (
            O => \N__30665\,
            I => \N__30662\
        );

    \I__5635\ : InMux
    port map (
            O => \N__30662\,
            I => \N__30658\
        );

    \I__5634\ : CascadeMux
    port map (
            O => \N__30661\,
            I => \N__30654\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__30658\,
            I => \N__30651\
        );

    \I__5632\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30648\
        );

    \I__5631\ : InMux
    port map (
            O => \N__30654\,
            I => \N__30645\
        );

    \I__5630\ : Span4Mux_h
    port map (
            O => \N__30651\,
            I => \N__30642\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__30648\,
            I => \N__30637\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__30645\,
            I => \N__30637\
        );

    \I__5627\ : Odrv4
    port map (
            O => \N__30642\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__30637\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__5625\ : InMux
    port map (
            O => \N__30632\,
            I => \bfn_12_22_0_\
        );

    \I__5624\ : InMux
    port map (
            O => \N__30629\,
            I => \N__30626\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__30626\,
            I => \N__30623\
        );

    \I__5622\ : Span4Mux_h
    port map (
            O => \N__30623\,
            I => \N__30619\
        );

    \I__5621\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30616\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__30619\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__30616\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__5618\ : InMux
    port map (
            O => \N__30611\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__5617\ : CascadeMux
    port map (
            O => \N__30608\,
            I => \N__30605\
        );

    \I__5616\ : InMux
    port map (
            O => \N__30605\,
            I => \N__30602\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__30602\,
            I => \N__30599\
        );

    \I__5614\ : Span4Mux_h
    port map (
            O => \N__30599\,
            I => \N__30595\
        );

    \I__5613\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30592\
        );

    \I__5612\ : Odrv4
    port map (
            O => \N__30595\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__30592\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__5610\ : InMux
    port map (
            O => \N__30587\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__5609\ : InMux
    port map (
            O => \N__30584\,
            I => \N__30581\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__30581\,
            I => \N__30577\
        );

    \I__5607\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30574\
        );

    \I__5606\ : Odrv4
    port map (
            O => \N__30577\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__30574\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__5604\ : InMux
    port map (
            O => \N__30569\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__5603\ : CascadeMux
    port map (
            O => \N__30566\,
            I => \N__30563\
        );

    \I__5602\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30560\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__30560\,
            I => \N__30556\
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__30559\,
            I => \N__30553\
        );

    \I__5599\ : Span4Mux_h
    port map (
            O => \N__30556\,
            I => \N__30550\
        );

    \I__5598\ : InMux
    port map (
            O => \N__30553\,
            I => \N__30547\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__30550\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__30547\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__5595\ : InMux
    port map (
            O => \N__30542\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__5594\ : CascadeMux
    port map (
            O => \N__30539\,
            I => \N__30536\
        );

    \I__5593\ : InMux
    port map (
            O => \N__30536\,
            I => \N__30533\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__30533\,
            I => \N__30530\
        );

    \I__5591\ : Span4Mux_v
    port map (
            O => \N__30530\,
            I => \N__30525\
        );

    \I__5590\ : InMux
    port map (
            O => \N__30529\,
            I => \N__30520\
        );

    \I__5589\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30520\
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__30525\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__30520\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__5586\ : InMux
    port map (
            O => \N__30515\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__5585\ : CascadeMux
    port map (
            O => \N__30512\,
            I => \N__30509\
        );

    \I__5584\ : InMux
    port map (
            O => \N__30509\,
            I => \N__30506\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__30506\,
            I => \N__30503\
        );

    \I__5582\ : Span4Mux_v
    port map (
            O => \N__30503\,
            I => \N__30498\
        );

    \I__5581\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30493\
        );

    \I__5580\ : InMux
    port map (
            O => \N__30501\,
            I => \N__30493\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__30498\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__30493\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5577\ : InMux
    port map (
            O => \N__30488\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__5576\ : CascadeMux
    port map (
            O => \N__30485\,
            I => \N__30482\
        );

    \I__5575\ : InMux
    port map (
            O => \N__30482\,
            I => \N__30479\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__30479\,
            I => \N__30476\
        );

    \I__5573\ : Span4Mux_v
    port map (
            O => \N__30476\,
            I => \N__30473\
        );

    \I__5572\ : Span4Mux_h
    port map (
            O => \N__30473\,
            I => \N__30467\
        );

    \I__5571\ : InMux
    port map (
            O => \N__30472\,
            I => \N__30464\
        );

    \I__5570\ : InMux
    port map (
            O => \N__30471\,
            I => \N__30461\
        );

    \I__5569\ : InMux
    port map (
            O => \N__30470\,
            I => \N__30458\
        );

    \I__5568\ : Odrv4
    port map (
            O => \N__30467\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__30464\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__30461\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__30458\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__5564\ : InMux
    port map (
            O => \N__30449\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__30446\,
            I => \N__30443\
        );

    \I__5562\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30440\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__30440\,
            I => \N__30436\
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__30439\,
            I => \N__30433\
        );

    \I__5559\ : Span4Mux_v
    port map (
            O => \N__30436\,
            I => \N__30430\
        );

    \I__5558\ : InMux
    port map (
            O => \N__30433\,
            I => \N__30427\
        );

    \I__5557\ : Odrv4
    port map (
            O => \N__30430\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__30427\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__5555\ : InMux
    port map (
            O => \N__30422\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__5554\ : CascadeMux
    port map (
            O => \N__30419\,
            I => \N__30416\
        );

    \I__5553\ : InMux
    port map (
            O => \N__30416\,
            I => \N__30413\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__30413\,
            I => \N__30410\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__30410\,
            I => \N__30406\
        );

    \I__5550\ : InMux
    port map (
            O => \N__30409\,
            I => \N__30403\
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__30406\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__30403\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__5547\ : InMux
    port map (
            O => \N__30398\,
            I => \bfn_12_21_0_\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__30395\,
            I => \N__30392\
        );

    \I__5545\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30389\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__30389\,
            I => \N__30386\
        );

    \I__5543\ : Span4Mux_v
    port map (
            O => \N__30386\,
            I => \N__30382\
        );

    \I__5542\ : InMux
    port map (
            O => \N__30385\,
            I => \N__30379\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__30382\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__30379\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__5539\ : InMux
    port map (
            O => \N__30374\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__30371\,
            I => \N__30368\
        );

    \I__5537\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30365\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__30365\,
            I => \N__30362\
        );

    \I__5535\ : Span4Mux_h
    port map (
            O => \N__30362\,
            I => \N__30358\
        );

    \I__5534\ : InMux
    port map (
            O => \N__30361\,
            I => \N__30355\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__30358\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__30355\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__5531\ : InMux
    port map (
            O => \N__30350\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__5530\ : CascadeMux
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__5529\ : InMux
    port map (
            O => \N__30344\,
            I => \N__30341\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__30341\,
            I => \N__30337\
        );

    \I__5527\ : InMux
    port map (
            O => \N__30340\,
            I => \N__30332\
        );

    \I__5526\ : Span4Mux_v
    port map (
            O => \N__30337\,
            I => \N__30329\
        );

    \I__5525\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30326\
        );

    \I__5524\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30323\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__30332\,
            I => \N__30320\
        );

    \I__5522\ : Span4Mux_h
    port map (
            O => \N__30329\,
            I => \N__30315\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__30326\,
            I => \N__30315\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__30323\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\
        );

    \I__5519\ : Odrv4
    port map (
            O => \N__30320\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__30315\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30308\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__5516\ : CascadeMux
    port map (
            O => \N__30305\,
            I => \N__30302\
        );

    \I__5515\ : InMux
    port map (
            O => \N__30302\,
            I => \N__30297\
        );

    \I__5514\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30294\
        );

    \I__5513\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30291\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__30297\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__30294\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__30291\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\
        );

    \I__5509\ : InMux
    port map (
            O => \N__30284\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__5508\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30277\
        );

    \I__5507\ : InMux
    port map (
            O => \N__30280\,
            I => \N__30274\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__30277\,
            I => \N__30271\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__30274\,
            I => \N__30267\
        );

    \I__5504\ : Span4Mux_h
    port map (
            O => \N__30271\,
            I => \N__30260\
        );

    \I__5503\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30257\
        );

    \I__5502\ : Span4Mux_h
    port map (
            O => \N__30267\,
            I => \N__30254\
        );

    \I__5501\ : InMux
    port map (
            O => \N__30266\,
            I => \N__30247\
        );

    \I__5500\ : InMux
    port map (
            O => \N__30265\,
            I => \N__30247\
        );

    \I__5499\ : InMux
    port map (
            O => \N__30264\,
            I => \N__30247\
        );

    \I__5498\ : InMux
    port map (
            O => \N__30263\,
            I => \N__30244\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__30260\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__30257\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__30254\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__30247\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__30244\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__5492\ : InMux
    port map (
            O => \N__30233\,
            I => \N__30228\
        );

    \I__5491\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30225\
        );

    \I__5490\ : CascadeMux
    port map (
            O => \N__30231\,
            I => \N__30222\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30228\,
            I => \N__30217\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__30225\,
            I => \N__30217\
        );

    \I__5487\ : InMux
    port map (
            O => \N__30222\,
            I => \N__30214\
        );

    \I__5486\ : Span4Mux_h
    port map (
            O => \N__30217\,
            I => \N__30211\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__30214\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__30211\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6\
        );

    \I__5483\ : InMux
    port map (
            O => \N__30206\,
            I => \N__30197\
        );

    \I__5482\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30194\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30204\,
            I => \N__30187\
        );

    \I__5480\ : InMux
    port map (
            O => \N__30203\,
            I => \N__30187\
        );

    \I__5479\ : InMux
    port map (
            O => \N__30202\,
            I => \N__30187\
        );

    \I__5478\ : InMux
    port map (
            O => \N__30201\,
            I => \N__30182\
        );

    \I__5477\ : InMux
    port map (
            O => \N__30200\,
            I => \N__30179\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__30197\,
            I => \N__30174\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__30194\,
            I => \N__30174\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__30187\,
            I => \N__30171\
        );

    \I__5473\ : InMux
    port map (
            O => \N__30186\,
            I => \N__30168\
        );

    \I__5472\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30165\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__30182\,
            I => \N__30162\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__30179\,
            I => \N__30157\
        );

    \I__5469\ : Span4Mux_v
    port map (
            O => \N__30174\,
            I => \N__30157\
        );

    \I__5468\ : Odrv12
    port map (
            O => \N__30171\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__30168\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__30165\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__5465\ : Odrv4
    port map (
            O => \N__30162\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__30157\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__30146\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_\
        );

    \I__5462\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30140\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__30140\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6\
        );

    \I__5460\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30134\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__30134\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6\
        );

    \I__5458\ : InMux
    port map (
            O => \N__30131\,
            I => \N__30125\
        );

    \I__5457\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30125\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__30125\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30122\,
            I => \N__30117\
        );

    \I__5454\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30112\
        );

    \I__5453\ : InMux
    port map (
            O => \N__30120\,
            I => \N__30112\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__30117\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__30112\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__30107\,
            I => \N__30104\
        );

    \I__5449\ : InMux
    port map (
            O => \N__30104\,
            I => \N__30101\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__30101\,
            I => \N__30098\
        );

    \I__5447\ : Span4Mux_v
    port map (
            O => \N__30098\,
            I => \N__30094\
        );

    \I__5446\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30091\
        );

    \I__5445\ : Odrv4
    port map (
            O => \N__30094\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__30091\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__5443\ : InMux
    port map (
            O => \N__30086\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__5442\ : CascadeMux
    port map (
            O => \N__30083\,
            I => \N__30080\
        );

    \I__5441\ : InMux
    port map (
            O => \N__30080\,
            I => \N__30077\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__30077\,
            I => \N__30074\
        );

    \I__5439\ : Span4Mux_h
    port map (
            O => \N__30074\,
            I => \N__30070\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30067\
        );

    \I__5437\ : Odrv4
    port map (
            O => \N__30070\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__30067\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__5435\ : InMux
    port map (
            O => \N__30062\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__5434\ : InMux
    port map (
            O => \N__30059\,
            I => \N__30052\
        );

    \I__5433\ : InMux
    port map (
            O => \N__30058\,
            I => \N__30052\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30049\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30052\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__30049\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\
        );

    \I__5429\ : InMux
    port map (
            O => \N__30044\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__5428\ : InMux
    port map (
            O => \N__30041\,
            I => \N__30038\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__30038\,
            I => \N__30035\
        );

    \I__5426\ : Span4Mux_h
    port map (
            O => \N__30035\,
            I => \N__30032\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__30032\,
            I => \phase_controller_inst1.stoper_hc.un6_running_17\
        );

    \I__5424\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30025\
        );

    \I__5423\ : InMux
    port map (
            O => \N__30028\,
            I => \N__30022\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__30025\,
            I => \N__30019\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__30022\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5420\ : Odrv12
    port map (
            O => \N__30019\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5419\ : CascadeMux
    port map (
            O => \N__30014\,
            I => \N__30011\
        );

    \I__5418\ : InMux
    port map (
            O => \N__30011\,
            I => \N__30008\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__30008\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30005\,
            I => \N__30002\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__30002\,
            I => \N__29999\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__29999\,
            I => \N__29996\
        );

    \I__5413\ : Odrv4
    port map (
            O => \N__29996\,
            I => \phase_controller_inst1.stoper_hc.un6_running_18\
        );

    \I__5412\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29989\
        );

    \I__5411\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29986\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__29989\,
            I => \N__29983\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__29986\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__5408\ : Odrv12
    port map (
            O => \N__29983\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__29978\,
            I => \N__29975\
        );

    \I__5406\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29972\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__29972\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__5404\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29966\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__29966\,
            I => \N__29963\
        );

    \I__5402\ : Span4Mux_v
    port map (
            O => \N__29963\,
            I => \N__29960\
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__29960\,
            I => \phase_controller_inst1.stoper_hc.un6_running_19\
        );

    \I__5400\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29953\
        );

    \I__5399\ : InMux
    port map (
            O => \N__29956\,
            I => \N__29950\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__29953\,
            I => \N__29947\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__29950\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__5396\ : Odrv4
    port map (
            O => \N__29947\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__5394\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29936\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__29936\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__5392\ : InMux
    port map (
            O => \N__29933\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_19\
        );

    \I__5391\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29926\
        );

    \I__5390\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29922\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__29926\,
            I => \N__29919\
        );

    \I__5388\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29916\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__29922\,
            I => \N__29913\
        );

    \I__5386\ : Span4Mux_h
    port map (
            O => \N__29919\,
            I => \N__29910\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__29916\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\
        );

    \I__5384\ : Odrv4
    port map (
            O => \N__29913\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\
        );

    \I__5383\ : Odrv4
    port map (
            O => \N__29910\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\
        );

    \I__5382\ : CascadeMux
    port map (
            O => \N__29903\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2_cascade_\
        );

    \I__5381\ : InMux
    port map (
            O => \N__29900\,
            I => \N__29897\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__29897\,
            I => \N__29893\
        );

    \I__5379\ : InMux
    port map (
            O => \N__29896\,
            I => \N__29890\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__29893\,
            I => \N__29887\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__29890\,
            I => \N__29884\
        );

    \I__5376\ : Odrv4
    port map (
            O => \N__29887\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\
        );

    \I__5375\ : Odrv4
    port map (
            O => \N__29884\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\
        );

    \I__5374\ : CascadeMux
    port map (
            O => \N__29879\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5_cascade_\
        );

    \I__5373\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29871\
        );

    \I__5372\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29865\
        );

    \I__5371\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29865\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__29871\,
            I => \N__29862\
        );

    \I__5369\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29859\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__29865\,
            I => \N__29856\
        );

    \I__5367\ : Span4Mux_h
    port map (
            O => \N__29862\,
            I => \N__29853\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__29859\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\
        );

    \I__5365\ : Odrv4
    port map (
            O => \N__29856\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\
        );

    \I__5364\ : Odrv4
    port map (
            O => \N__29853\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\
        );

    \I__5363\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29843\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__29843\,
            I => \N__29840\
        );

    \I__5361\ : Span4Mux_h
    port map (
            O => \N__29840\,
            I => \N__29837\
        );

    \I__5360\ : Odrv4
    port map (
            O => \N__29837\,
            I => \phase_controller_inst1.stoper_hc.un6_running_9\
        );

    \I__5359\ : InMux
    port map (
            O => \N__29834\,
            I => \N__29830\
        );

    \I__5358\ : InMux
    port map (
            O => \N__29833\,
            I => \N__29827\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__29830\,
            I => \N__29824\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__29827\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5355\ : Odrv12
    port map (
            O => \N__29824\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__29819\,
            I => \N__29816\
        );

    \I__5353\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29813\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__29813\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__5351\ : CascadeMux
    port map (
            O => \N__29810\,
            I => \N__29807\
        );

    \I__5350\ : InMux
    port map (
            O => \N__29807\,
            I => \N__29804\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__29804\,
            I => \N__29801\
        );

    \I__5348\ : Span4Mux_h
    port map (
            O => \N__29801\,
            I => \N__29798\
        );

    \I__5347\ : Odrv4
    port map (
            O => \N__29798\,
            I => \phase_controller_inst1.stoper_hc.un6_running_10\
        );

    \I__5346\ : InMux
    port map (
            O => \N__29795\,
            I => \N__29791\
        );

    \I__5345\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29788\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__29791\,
            I => \N__29785\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__29788\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__5342\ : Odrv12
    port map (
            O => \N__29785\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__5341\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29777\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__29777\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__5339\ : CascadeMux
    port map (
            O => \N__29774\,
            I => \N__29771\
        );

    \I__5338\ : InMux
    port map (
            O => \N__29771\,
            I => \N__29768\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__29768\,
            I => \phase_controller_inst1.stoper_hc.un6_running_11\
        );

    \I__5336\ : InMux
    port map (
            O => \N__29765\,
            I => \N__29761\
        );

    \I__5335\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29758\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__29761\,
            I => \N__29755\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__29758\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__5332\ : Odrv4
    port map (
            O => \N__29755\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__5331\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29747\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__29747\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__5329\ : CascadeMux
    port map (
            O => \N__29744\,
            I => \N__29741\
        );

    \I__5328\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29738\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__29738\,
            I => \phase_controller_inst1.stoper_hc.un6_running_12\
        );

    \I__5326\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29731\
        );

    \I__5325\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29728\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__29731\,
            I => \N__29725\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__29728\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__29725\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5321\ : InMux
    port map (
            O => \N__29720\,
            I => \N__29717\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__29717\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__5319\ : CascadeMux
    port map (
            O => \N__29714\,
            I => \N__29711\
        );

    \I__5318\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29708\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__29708\,
            I => \phase_controller_inst1.stoper_hc.un6_running_13\
        );

    \I__5316\ : InMux
    port map (
            O => \N__29705\,
            I => \N__29701\
        );

    \I__5315\ : InMux
    port map (
            O => \N__29704\,
            I => \N__29698\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__29701\,
            I => \N__29695\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__29698\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5312\ : Odrv4
    port map (
            O => \N__29695\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5311\ : InMux
    port map (
            O => \N__29690\,
            I => \N__29687\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__29687\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__5309\ : InMux
    port map (
            O => \N__29684\,
            I => \N__29681\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__29681\,
            I => \N__29678\
        );

    \I__5307\ : Span12Mux_h
    port map (
            O => \N__29678\,
            I => \N__29675\
        );

    \I__5306\ : Odrv12
    port map (
            O => \N__29675\,
            I => \phase_controller_inst1.stoper_hc.un6_running_14\
        );

    \I__5305\ : InMux
    port map (
            O => \N__29672\,
            I => \N__29668\
        );

    \I__5304\ : InMux
    port map (
            O => \N__29671\,
            I => \N__29665\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__29668\,
            I => \N__29662\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__29665\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5301\ : Odrv4
    port map (
            O => \N__29662\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5300\ : CascadeMux
    port map (
            O => \N__29657\,
            I => \N__29654\
        );

    \I__5299\ : InMux
    port map (
            O => \N__29654\,
            I => \N__29651\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__29651\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__5297\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29644\
        );

    \I__5296\ : InMux
    port map (
            O => \N__29647\,
            I => \N__29641\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__29644\,
            I => \N__29638\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__29641\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__29638\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__5292\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29630\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__29630\,
            I => \phase_controller_inst1.stoper_hc.un6_running_15\
        );

    \I__5290\ : CascadeMux
    port map (
            O => \N__29627\,
            I => \N__29624\
        );

    \I__5289\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29621\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__29621\,
            I => \N__29618\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__29618\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__5286\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29612\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__29612\,
            I => \N__29609\
        );

    \I__5284\ : Span12Mux_v
    port map (
            O => \N__29609\,
            I => \N__29606\
        );

    \I__5283\ : Odrv12
    port map (
            O => \N__29606\,
            I => \phase_controller_inst1.stoper_hc.un6_running_16\
        );

    \I__5282\ : InMux
    port map (
            O => \N__29603\,
            I => \N__29599\
        );

    \I__5281\ : InMux
    port map (
            O => \N__29602\,
            I => \N__29596\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__29599\,
            I => \N__29593\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__29596\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__29593\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5277\ : CascadeMux
    port map (
            O => \N__29588\,
            I => \N__29585\
        );

    \I__5276\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29582\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__29582\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__5274\ : InMux
    port map (
            O => \N__29579\,
            I => \N__29576\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__29576\,
            I => \N__29573\
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__29573\,
            I => \phase_controller_inst1.stoper_hc.un6_running_2\
        );

    \I__5271\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29567\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__29567\,
            I => \N__29563\
        );

    \I__5269\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29560\
        );

    \I__5268\ : Span4Mux_v
    port map (
            O => \N__29563\,
            I => \N__29557\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__29560\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__5266\ : Odrv4
    port map (
            O => \N__29557\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__5265\ : CascadeMux
    port map (
            O => \N__29552\,
            I => \N__29549\
        );

    \I__5264\ : InMux
    port map (
            O => \N__29549\,
            I => \N__29546\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__29546\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__5262\ : InMux
    port map (
            O => \N__29543\,
            I => \N__29540\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__29540\,
            I => \phase_controller_inst1.stoper_hc.un6_running_3\
        );

    \I__5260\ : CascadeMux
    port map (
            O => \N__29537\,
            I => \N__29533\
        );

    \I__5259\ : InMux
    port map (
            O => \N__29536\,
            I => \N__29530\
        );

    \I__5258\ : InMux
    port map (
            O => \N__29533\,
            I => \N__29527\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__29530\,
            I => \N__29524\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__29527\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__29524\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__5254\ : CascadeMux
    port map (
            O => \N__29519\,
            I => \N__29516\
        );

    \I__5253\ : InMux
    port map (
            O => \N__29516\,
            I => \N__29513\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__29513\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__5251\ : InMux
    port map (
            O => \N__29510\,
            I => \N__29506\
        );

    \I__5250\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29503\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__29506\,
            I => \N__29500\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__29503\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__29500\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__5246\ : InMux
    port map (
            O => \N__29495\,
            I => \N__29492\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__29492\,
            I => \N__29489\
        );

    \I__5244\ : Odrv4
    port map (
            O => \N__29489\,
            I => \phase_controller_inst1.stoper_hc.un6_running_4\
        );

    \I__5243\ : CascadeMux
    port map (
            O => \N__29486\,
            I => \N__29483\
        );

    \I__5242\ : InMux
    port map (
            O => \N__29483\,
            I => \N__29480\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__29480\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__5240\ : InMux
    port map (
            O => \N__29477\,
            I => \N__29474\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__29474\,
            I => \N__29471\
        );

    \I__5238\ : Odrv4
    port map (
            O => \N__29471\,
            I => \phase_controller_inst1.stoper_hc.un6_running_5\
        );

    \I__5237\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29464\
        );

    \I__5236\ : InMux
    port map (
            O => \N__29467\,
            I => \N__29461\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__29464\,
            I => \N__29458\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__29461\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5233\ : Odrv4
    port map (
            O => \N__29458\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5232\ : CascadeMux
    port map (
            O => \N__29453\,
            I => \N__29450\
        );

    \I__5231\ : InMux
    port map (
            O => \N__29450\,
            I => \N__29447\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__29447\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__5229\ : InMux
    port map (
            O => \N__29444\,
            I => \N__29441\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__29441\,
            I => \N__29438\
        );

    \I__5227\ : Odrv4
    port map (
            O => \N__29438\,
            I => \phase_controller_inst1.stoper_hc.un6_running_6\
        );

    \I__5226\ : InMux
    port map (
            O => \N__29435\,
            I => \N__29431\
        );

    \I__5225\ : InMux
    port map (
            O => \N__29434\,
            I => \N__29428\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__29431\,
            I => \N__29425\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__29428\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5222\ : Odrv4
    port map (
            O => \N__29425\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5221\ : CascadeMux
    port map (
            O => \N__29420\,
            I => \N__29417\
        );

    \I__5220\ : InMux
    port map (
            O => \N__29417\,
            I => \N__29414\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__29414\,
            I => \N__29411\
        );

    \I__5218\ : Odrv4
    port map (
            O => \N__29411\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__5217\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29404\
        );

    \I__5216\ : InMux
    port map (
            O => \N__29407\,
            I => \N__29401\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__29404\,
            I => \N__29398\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__29401\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__29398\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__29393\,
            I => \N__29390\
        );

    \I__5211\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29387\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__29387\,
            I => \phase_controller_inst1.stoper_hc.un6_running_7\
        );

    \I__5209\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29381\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__29381\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__5207\ : CascadeMux
    port map (
            O => \N__29378\,
            I => \N__29375\
        );

    \I__5206\ : InMux
    port map (
            O => \N__29375\,
            I => \N__29372\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__29372\,
            I => \phase_controller_inst1.stoper_hc.un6_running_8\
        );

    \I__5204\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29365\
        );

    \I__5203\ : InMux
    port map (
            O => \N__29368\,
            I => \N__29362\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__29365\,
            I => \N__29359\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__29362\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5200\ : Odrv4
    port map (
            O => \N__29359\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5199\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29351\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__29351\,
            I => \N__29348\
        );

    \I__5197\ : Odrv4
    port map (
            O => \N__29348\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29345\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__5195\ : InMux
    port map (
            O => \N__29342\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__5194\ : InMux
    port map (
            O => \N__29339\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__5193\ : InMux
    port map (
            O => \N__29336\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__5192\ : InMux
    port map (
            O => \N__29333\,
            I => \bfn_12_15_0_\
        );

    \I__5191\ : InMux
    port map (
            O => \N__29330\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__5190\ : InMux
    port map (
            O => \N__29327\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__5189\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29321\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__29321\,
            I => \N__29317\
        );

    \I__5187\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29314\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__29317\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__29314\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__5184\ : CEMux
    port map (
            O => \N__29309\,
            I => \N__29305\
        );

    \I__5183\ : CEMux
    port map (
            O => \N__29308\,
            I => \N__29301\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__29305\,
            I => \N__29294\
        );

    \I__5181\ : CEMux
    port map (
            O => \N__29304\,
            I => \N__29291\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__29301\,
            I => \N__29288\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29300\,
            I => \N__29268\
        );

    \I__5178\ : InMux
    port map (
            O => \N__29299\,
            I => \N__29268\
        );

    \I__5177\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29263\
        );

    \I__5176\ : InMux
    port map (
            O => \N__29297\,
            I => \N__29263\
        );

    \I__5175\ : Span4Mux_v
    port map (
            O => \N__29294\,
            I => \N__29258\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__29291\,
            I => \N__29258\
        );

    \I__5173\ : Span4Mux_v
    port map (
            O => \N__29288\,
            I => \N__29255\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29287\,
            I => \N__29246\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29286\,
            I => \N__29246\
        );

    \I__5170\ : InMux
    port map (
            O => \N__29285\,
            I => \N__29246\
        );

    \I__5169\ : InMux
    port map (
            O => \N__29284\,
            I => \N__29246\
        );

    \I__5168\ : InMux
    port map (
            O => \N__29283\,
            I => \N__29237\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29237\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29281\,
            I => \N__29237\
        );

    \I__5165\ : InMux
    port map (
            O => \N__29280\,
            I => \N__29237\
        );

    \I__5164\ : InMux
    port map (
            O => \N__29279\,
            I => \N__29230\
        );

    \I__5163\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29230\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29230\
        );

    \I__5161\ : InMux
    port map (
            O => \N__29276\,
            I => \N__29221\
        );

    \I__5160\ : InMux
    port map (
            O => \N__29275\,
            I => \N__29221\
        );

    \I__5159\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29221\
        );

    \I__5158\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29221\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__29268\,
            I => \N__29214\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__29263\,
            I => \N__29214\
        );

    \I__5155\ : Span4Mux_h
    port map (
            O => \N__29258\,
            I => \N__29214\
        );

    \I__5154\ : Span4Mux_h
    port map (
            O => \N__29255\,
            I => \N__29211\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__29246\,
            I => \N__29208\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__29237\,
            I => \N__29199\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__29230\,
            I => \N__29199\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__29221\,
            I => \N__29199\
        );

    \I__5149\ : Span4Mux_v
    port map (
            O => \N__29214\,
            I => \N__29199\
        );

    \I__5148\ : Span4Mux_v
    port map (
            O => \N__29211\,
            I => \N__29196\
        );

    \I__5147\ : Span4Mux_v
    port map (
            O => \N__29208\,
            I => \N__29191\
        );

    \I__5146\ : Span4Mux_v
    port map (
            O => \N__29199\,
            I => \N__29191\
        );

    \I__5145\ : Span4Mux_v
    port map (
            O => \N__29196\,
            I => \N__29188\
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__29191\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__5143\ : Odrv4
    port map (
            O => \N__29188\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__5142\ : InMux
    port map (
            O => \N__29183\,
            I => \N__29180\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29180\,
            I => \N__29177\
        );

    \I__5140\ : Span4Mux_v
    port map (
            O => \N__29177\,
            I => \N__29174\
        );

    \I__5139\ : Span4Mux_h
    port map (
            O => \N__29174\,
            I => \N__29171\
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__29171\,
            I => \phase_controller_inst1.stoper_hc.un6_running_1\
        );

    \I__5137\ : CascadeMux
    port map (
            O => \N__29168\,
            I => \N__29164\
        );

    \I__5136\ : InMux
    port map (
            O => \N__29167\,
            I => \N__29161\
        );

    \I__5135\ : InMux
    port map (
            O => \N__29164\,
            I => \N__29157\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__29161\,
            I => \N__29154\
        );

    \I__5133\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29151\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__29157\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__29154\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__29151\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5129\ : CascadeMux
    port map (
            O => \N__29144\,
            I => \N__29141\
        );

    \I__5128\ : InMux
    port map (
            O => \N__29141\,
            I => \N__29138\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__29138\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__5126\ : InMux
    port map (
            O => \N__29135\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__5125\ : InMux
    port map (
            O => \N__29132\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__5124\ : InMux
    port map (
            O => \N__29129\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__5123\ : InMux
    port map (
            O => \N__29126\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__5122\ : InMux
    port map (
            O => \N__29123\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29120\,
            I => \bfn_12_14_0_\
        );

    \I__5120\ : InMux
    port map (
            O => \N__29117\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__5119\ : InMux
    port map (
            O => \N__29114\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29111\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__5117\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29105\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__29105\,
            I => \N__29101\
        );

    \I__5115\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29098\
        );

    \I__5114\ : Span4Mux_v
    port map (
            O => \N__29101\,
            I => \N__29092\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29092\
        );

    \I__5112\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29089\
        );

    \I__5111\ : Odrv4
    port map (
            O => \N__29092\,
            I => \il_min_comp1_D2\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__29089\,
            I => \il_min_comp1_D2\
        );

    \I__5109\ : InMux
    port map (
            O => \N__29084\,
            I => \N__29080\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29083\,
            I => \N__29077\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__29080\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__29077\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__5105\ : InMux
    port map (
            O => \N__29072\,
            I => \N__29068\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29065\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29059\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__29065\,
            I => \N__29059\
        );

    \I__5101\ : InMux
    port map (
            O => \N__29064\,
            I => \N__29056\
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__29059\,
            I => \il_max_comp1_D2\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__29056\,
            I => \il_max_comp1_D2\
        );

    \I__5098\ : InMux
    port map (
            O => \N__29051\,
            I => \N__29045\
        );

    \I__5097\ : InMux
    port map (
            O => \N__29050\,
            I => \N__29045\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__29045\,
            I => \phase_controller_inst1.N_56\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__29042\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__5094\ : CascadeMux
    port map (
            O => \N__29039\,
            I => \N__29036\
        );

    \I__5093\ : InMux
    port map (
            O => \N__29036\,
            I => \N__29033\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__29033\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__5091\ : InMux
    port map (
            O => \N__29030\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__5090\ : InMux
    port map (
            O => \N__29027\,
            I => \N__29024\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__29024\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3DZ0Z41\
        );

    \I__5088\ : InMux
    port map (
            O => \N__29021\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__5087\ : InMux
    port map (
            O => \N__29018\,
            I => \N__29015\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__29015\,
            I => \N__29012\
        );

    \I__5085\ : Span4Mux_v
    port map (
            O => \N__29012\,
            I => \N__29009\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__29009\,
            I => \il_max_comp1_D1\
        );

    \I__5083\ : InMux
    port map (
            O => \N__29006\,
            I => \N__29003\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__29003\,
            I => \N__29000\
        );

    \I__5081\ : Odrv12
    port map (
            O => \N__29000\,
            I => \il_min_comp2_D1\
        );

    \I__5080\ : InMux
    port map (
            O => \N__28997\,
            I => \N__28994\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__28994\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__5078\ : InMux
    port map (
            O => \N__28991\,
            I => \N__28988\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__28988\,
            I => \phase_controller_inst1.N_55\
        );

    \I__5076\ : InMux
    port map (
            O => \N__28985\,
            I => \N__28978\
        );

    \I__5075\ : InMux
    port map (
            O => \N__28984\,
            I => \N__28978\
        );

    \I__5074\ : InMux
    port map (
            O => \N__28983\,
            I => \N__28975\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__28978\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__28975\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5071\ : CascadeMux
    port map (
            O => \N__28970\,
            I => \N__28966\
        );

    \I__5070\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28959\
        );

    \I__5069\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28959\
        );

    \I__5068\ : InMux
    port map (
            O => \N__28965\,
            I => \N__28956\
        );

    \I__5067\ : InMux
    port map (
            O => \N__28964\,
            I => \N__28953\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__28959\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__28956\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__28953\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5063\ : InMux
    port map (
            O => \N__28946\,
            I => \N__28943\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__28943\,
            I => \N__28940\
        );

    \I__5061\ : Span4Mux_h
    port map (
            O => \N__28940\,
            I => \N__28937\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__28937\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__5059\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28931\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__28931\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5\
        );

    \I__5057\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28921\
        );

    \I__5056\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28921\
        );

    \I__5055\ : InMux
    port map (
            O => \N__28926\,
            I => \N__28918\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__28921\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__28918\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO\
        );

    \I__5052\ : InMux
    port map (
            O => \N__28913\,
            I => \N__28909\
        );

    \I__5051\ : InMux
    port map (
            O => \N__28912\,
            I => \N__28906\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__28909\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__28906\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__5048\ : CascadeMux
    port map (
            O => \N__28901\,
            I => \N__28898\
        );

    \I__5047\ : InMux
    port map (
            O => \N__28898\,
            I => \N__28893\
        );

    \I__5046\ : InMux
    port map (
            O => \N__28897\,
            I => \N__28890\
        );

    \I__5045\ : InMux
    port map (
            O => \N__28896\,
            I => \N__28887\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__28893\,
            I => \N__28884\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__28890\,
            I => \N__28881\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__28887\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__28884\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5040\ : Odrv4
    port map (
            O => \N__28881\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5039\ : CEMux
    port map (
            O => \N__28874\,
            I => \N__28863\
        );

    \I__5038\ : CEMux
    port map (
            O => \N__28873\,
            I => \N__28859\
        );

    \I__5037\ : CEMux
    port map (
            O => \N__28872\,
            I => \N__28856\
        );

    \I__5036\ : CEMux
    port map (
            O => \N__28871\,
            I => \N__28853\
        );

    \I__5035\ : InMux
    port map (
            O => \N__28870\,
            I => \N__28844\
        );

    \I__5034\ : InMux
    port map (
            O => \N__28869\,
            I => \N__28844\
        );

    \I__5033\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28844\
        );

    \I__5032\ : InMux
    port map (
            O => \N__28867\,
            I => \N__28844\
        );

    \I__5031\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28841\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__28863\,
            I => \N__28838\
        );

    \I__5029\ : CEMux
    port map (
            O => \N__28862\,
            I => \N__28835\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__28859\,
            I => \N__28830\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__28856\,
            I => \N__28830\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__28853\,
            I => \N__28825\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__28844\,
            I => \N__28808\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__28841\,
            I => \N__28808\
        );

    \I__5023\ : Sp12to4
    port map (
            O => \N__28838\,
            I => \N__28805\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__28835\,
            I => \N__28802\
        );

    \I__5021\ : Span4Mux_h
    port map (
            O => \N__28830\,
            I => \N__28799\
        );

    \I__5020\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28794\
        );

    \I__5019\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28794\
        );

    \I__5018\ : Span4Mux_h
    port map (
            O => \N__28825\,
            I => \N__28791\
        );

    \I__5017\ : InMux
    port map (
            O => \N__28824\,
            I => \N__28784\
        );

    \I__5016\ : InMux
    port map (
            O => \N__28823\,
            I => \N__28784\
        );

    \I__5015\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28784\
        );

    \I__5014\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28781\
        );

    \I__5013\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28772\
        );

    \I__5012\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28772\
        );

    \I__5011\ : InMux
    port map (
            O => \N__28818\,
            I => \N__28772\
        );

    \I__5010\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28772\
        );

    \I__5009\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28763\
        );

    \I__5008\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28763\
        );

    \I__5007\ : InMux
    port map (
            O => \N__28814\,
            I => \N__28763\
        );

    \I__5006\ : InMux
    port map (
            O => \N__28813\,
            I => \N__28763\
        );

    \I__5005\ : Span12Mux_s6_v
    port map (
            O => \N__28808\,
            I => \N__28758\
        );

    \I__5004\ : Span12Mux_v
    port map (
            O => \N__28805\,
            I => \N__28758\
        );

    \I__5003\ : Span4Mux_h
    port map (
            O => \N__28802\,
            I => \N__28753\
        );

    \I__5002\ : Span4Mux_v
    port map (
            O => \N__28799\,
            I => \N__28753\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__28794\,
            I => \N__28748\
        );

    \I__5000\ : Span4Mux_v
    port map (
            O => \N__28791\,
            I => \N__28748\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__28784\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__28781\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__28772\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__28763\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4995\ : Odrv12
    port map (
            O => \N__28758\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__28753\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4993\ : Odrv4
    port map (
            O => \N__28748\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4992\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28729\
        );

    \I__4991\ : InMux
    port map (
            O => \N__28732\,
            I => \N__28726\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__28729\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__28726\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__4988\ : CascadeMux
    port map (
            O => \N__28721\,
            I => \N__28717\
        );

    \I__4987\ : CascadeMux
    port map (
            O => \N__28720\,
            I => \N__28714\
        );

    \I__4986\ : InMux
    port map (
            O => \N__28717\,
            I => \N__28708\
        );

    \I__4985\ : InMux
    port map (
            O => \N__28714\,
            I => \N__28703\
        );

    \I__4984\ : InMux
    port map (
            O => \N__28713\,
            I => \N__28703\
        );

    \I__4983\ : InMux
    port map (
            O => \N__28712\,
            I => \N__28698\
        );

    \I__4982\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28698\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__28708\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__28703\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__28698\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__4978\ : InMux
    port map (
            O => \N__28691\,
            I => \N__28686\
        );

    \I__4977\ : InMux
    port map (
            O => \N__28690\,
            I => \N__28682\
        );

    \I__4976\ : InMux
    port map (
            O => \N__28689\,
            I => \N__28679\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__28686\,
            I => \N__28676\
        );

    \I__4974\ : InMux
    port map (
            O => \N__28685\,
            I => \N__28673\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__28682\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__28679\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4971\ : Odrv4
    port map (
            O => \N__28676\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__28673\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4969\ : IoInMux
    port map (
            O => \N__28664\,
            I => \N__28661\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__28661\,
            I => \N__28658\
        );

    \I__4967\ : Span4Mux_s1_v
    port map (
            O => \N__28658\,
            I => \N__28655\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__28655\,
            I => s4_phy_c
        );

    \I__4965\ : CascadeMux
    port map (
            O => \N__28652\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_\
        );

    \I__4964\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28646\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__28646\,
            I => \N__28640\
        );

    \I__4962\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28637\
        );

    \I__4961\ : InMux
    port map (
            O => \N__28644\,
            I => \N__28634\
        );

    \I__4960\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28631\
        );

    \I__4959\ : Span4Mux_h
    port map (
            O => \N__28640\,
            I => \N__28628\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__28637\,
            I => \N__28623\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__28634\,
            I => \N__28623\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__28631\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__28628\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3\
        );

    \I__4954\ : Odrv4
    port map (
            O => \N__28623\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3\
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__28616\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3_cascade_\
        );

    \I__4952\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28610\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__28610\,
            I => \N__28607\
        );

    \I__4950\ : Odrv4
    port map (
            O => \N__28607\,
            I => \phase_controller_inst1.stoper_hc.N_283\
        );

    \I__4949\ : InMux
    port map (
            O => \N__28604\,
            I => \N__28598\
        );

    \I__4948\ : InMux
    port map (
            O => \N__28603\,
            I => \N__28598\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__28598\,
            I => \N__28595\
        );

    \I__4946\ : Span4Mux_v
    port map (
            O => \N__28595\,
            I => \N__28591\
        );

    \I__4945\ : InMux
    port map (
            O => \N__28594\,
            I => \N__28588\
        );

    \I__4944\ : Odrv4
    port map (
            O => \N__28591\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__28588\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\
        );

    \I__4942\ : CascadeMux
    port map (
            O => \N__28583\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_\
        );

    \I__4941\ : InMux
    port map (
            O => \N__28580\,
            I => \N__28577\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__28577\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15\
        );

    \I__4939\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28571\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__28571\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10\
        );

    \I__4937\ : CascadeMux
    port map (
            O => \N__28568\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_\
        );

    \I__4936\ : CascadeMux
    port map (
            O => \N__28565\,
            I => \N__28561\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__28564\,
            I => \N__28558\
        );

    \I__4934\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28553\
        );

    \I__4933\ : InMux
    port map (
            O => \N__28558\,
            I => \N__28553\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__28553\,
            I => \N__28549\
        );

    \I__4931\ : InMux
    port map (
            O => \N__28552\,
            I => \N__28546\
        );

    \I__4930\ : Span4Mux_h
    port map (
            O => \N__28549\,
            I => \N__28543\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__28546\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__28543\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\
        );

    \I__4927\ : InMux
    port map (
            O => \N__28538\,
            I => \N__28535\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__28535\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4\
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__28532\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_\
        );

    \I__4924\ : InMux
    port map (
            O => \N__28529\,
            I => \N__28526\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__28526\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31\
        );

    \I__4922\ : CascadeMux
    port map (
            O => \N__28523\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i_cascade_\
        );

    \I__4921\ : InMux
    port map (
            O => \N__28520\,
            I => \N__28516\
        );

    \I__4920\ : InMux
    port map (
            O => \N__28519\,
            I => \N__28513\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__28516\,
            I => \elapsed_time_ns_1_RNIS5ND11_0_24\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__28513\,
            I => \elapsed_time_ns_1_RNIS5ND11_0_24\
        );

    \I__4917\ : InMux
    port map (
            O => \N__28508\,
            I => \N__28504\
        );

    \I__4916\ : InMux
    port map (
            O => \N__28507\,
            I => \N__28501\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__28504\,
            I => \elapsed_time_ns_1_RNIT6ND11_0_25\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__28501\,
            I => \elapsed_time_ns_1_RNIT6ND11_0_25\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__28496\,
            I => \N__28491\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__28495\,
            I => \N__28486\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__28494\,
            I => \N__28482\
        );

    \I__4910\ : InMux
    port map (
            O => \N__28491\,
            I => \N__28477\
        );

    \I__4909\ : InMux
    port map (
            O => \N__28490\,
            I => \N__28474\
        );

    \I__4908\ : InMux
    port map (
            O => \N__28489\,
            I => \N__28471\
        );

    \I__4907\ : InMux
    port map (
            O => \N__28486\,
            I => \N__28468\
        );

    \I__4906\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28465\
        );

    \I__4905\ : InMux
    port map (
            O => \N__28482\,
            I => \N__28462\
        );

    \I__4904\ : InMux
    port map (
            O => \N__28481\,
            I => \N__28458\
        );

    \I__4903\ : InMux
    port map (
            O => \N__28480\,
            I => \N__28455\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__28477\,
            I => \N__28452\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__28474\,
            I => \N__28447\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__28471\,
            I => \N__28447\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__28468\,
            I => \N__28444\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__28465\,
            I => \N__28439\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__28462\,
            I => \N__28439\
        );

    \I__4896\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28436\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__28458\,
            I => \N__28433\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__28455\,
            I => \N__28426\
        );

    \I__4893\ : Span4Mux_h
    port map (
            O => \N__28452\,
            I => \N__28426\
        );

    \I__4892\ : Span4Mux_h
    port map (
            O => \N__28447\,
            I => \N__28426\
        );

    \I__4891\ : Span4Mux_v
    port map (
            O => \N__28444\,
            I => \N__28421\
        );

    \I__4890\ : Span4Mux_h
    port map (
            O => \N__28439\,
            I => \N__28421\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__28436\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__4888\ : Odrv12
    port map (
            O => \N__28433\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__28426\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__28421\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__4885\ : CascadeMux
    port map (
            O => \N__28412\,
            I => \N__28408\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__28411\,
            I => \N__28405\
        );

    \I__4883\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28402\
        );

    \I__4882\ : InMux
    port map (
            O => \N__28405\,
            I => \N__28399\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__28402\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__28399\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16\
        );

    \I__4879\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28390\
        );

    \I__4878\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28387\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__28390\,
            I => \elapsed_time_ns_1_RNIQ3ND11_0_22\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__28387\,
            I => \elapsed_time_ns_1_RNIQ3ND11_0_22\
        );

    \I__4875\ : CascadeMux
    port map (
            O => \N__28382\,
            I => \N__28379\
        );

    \I__4874\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28375\
        );

    \I__4873\ : InMux
    port map (
            O => \N__28378\,
            I => \N__28372\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__28375\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__28372\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__28367\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_\
        );

    \I__4869\ : CascadeMux
    port map (
            O => \N__28364\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_\
        );

    \I__4868\ : CascadeMux
    port map (
            O => \N__28361\,
            I => \N__28358\
        );

    \I__4867\ : InMux
    port map (
            O => \N__28358\,
            I => \N__28355\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__28355\,
            I => \N__28351\
        );

    \I__4865\ : InMux
    port map (
            O => \N__28354\,
            I => \N__28348\
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__28351\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__28348\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__28343\,
            I => \N__28340\
        );

    \I__4861\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28334\
        );

    \I__4860\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28331\
        );

    \I__4859\ : InMux
    port map (
            O => \N__28338\,
            I => \N__28328\
        );

    \I__4858\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28325\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__28334\,
            I => \N__28320\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__28331\,
            I => \N__28320\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__28328\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__28325\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4\
        );

    \I__4853\ : Odrv4
    port map (
            O => \N__28320\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4\
        );

    \I__4852\ : InMux
    port map (
            O => \N__28313\,
            I => \N__28299\
        );

    \I__4851\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28299\
        );

    \I__4850\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28299\
        );

    \I__4849\ : CascadeMux
    port map (
            O => \N__28310\,
            I => \N__28295\
        );

    \I__4848\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28281\
        );

    \I__4847\ : InMux
    port map (
            O => \N__28308\,
            I => \N__28281\
        );

    \I__4846\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28281\
        );

    \I__4845\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28281\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__28299\,
            I => \N__28278\
        );

    \I__4843\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28273\
        );

    \I__4842\ : InMux
    port map (
            O => \N__28295\,
            I => \N__28273\
        );

    \I__4841\ : InMux
    port map (
            O => \N__28294\,
            I => \N__28262\
        );

    \I__4840\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28262\
        );

    \I__4839\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28262\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28262\
        );

    \I__4837\ : InMux
    port map (
            O => \N__28290\,
            I => \N__28262\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__28281\,
            I => \N__28259\
        );

    \I__4835\ : Span4Mux_h
    port map (
            O => \N__28278\,
            I => \N__28256\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__28273\,
            I => \phase_controller_inst1.stoper_hc.N_325\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__28262\,
            I => \phase_controller_inst1.stoper_hc.N_325\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__28259\,
            I => \phase_controller_inst1.stoper_hc.N_325\
        );

    \I__4831\ : Odrv4
    port map (
            O => \N__28256\,
            I => \phase_controller_inst1.stoper_hc.N_325\
        );

    \I__4830\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28215\
        );

    \I__4829\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28215\
        );

    \I__4828\ : InMux
    port map (
            O => \N__28245\,
            I => \N__28215\
        );

    \I__4827\ : InMux
    port map (
            O => \N__28244\,
            I => \N__28215\
        );

    \I__4826\ : InMux
    port map (
            O => \N__28243\,
            I => \N__28215\
        );

    \I__4825\ : InMux
    port map (
            O => \N__28242\,
            I => \N__28212\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28201\
        );

    \I__4823\ : InMux
    port map (
            O => \N__28240\,
            I => \N__28201\
        );

    \I__4822\ : InMux
    port map (
            O => \N__28239\,
            I => \N__28201\
        );

    \I__4821\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28201\
        );

    \I__4820\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28201\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28236\,
            I => \N__28186\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28235\,
            I => \N__28186\
        );

    \I__4817\ : InMux
    port map (
            O => \N__28234\,
            I => \N__28186\
        );

    \I__4816\ : InMux
    port map (
            O => \N__28233\,
            I => \N__28186\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28232\,
            I => \N__28186\
        );

    \I__4814\ : InMux
    port map (
            O => \N__28231\,
            I => \N__28186\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28230\,
            I => \N__28186\
        );

    \I__4812\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28177\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28228\,
            I => \N__28177\
        );

    \I__4810\ : InMux
    port map (
            O => \N__28227\,
            I => \N__28177\
        );

    \I__4809\ : InMux
    port map (
            O => \N__28226\,
            I => \N__28177\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__28215\,
            I => \N__28160\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__28212\,
            I => \N__28157\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__28201\,
            I => \N__28150\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__28186\,
            I => \N__28150\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__28177\,
            I => \N__28150\
        );

    \I__4803\ : InMux
    port map (
            O => \N__28176\,
            I => \N__28147\
        );

    \I__4802\ : InMux
    port map (
            O => \N__28175\,
            I => \N__28140\
        );

    \I__4801\ : InMux
    port map (
            O => \N__28174\,
            I => \N__28140\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28140\
        );

    \I__4799\ : InMux
    port map (
            O => \N__28172\,
            I => \N__28127\
        );

    \I__4798\ : InMux
    port map (
            O => \N__28171\,
            I => \N__28127\
        );

    \I__4797\ : InMux
    port map (
            O => \N__28170\,
            I => \N__28127\
        );

    \I__4796\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28127\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28168\,
            I => \N__28127\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28127\
        );

    \I__4793\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28118\
        );

    \I__4792\ : InMux
    port map (
            O => \N__28165\,
            I => \N__28118\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28118\
        );

    \I__4790\ : InMux
    port map (
            O => \N__28163\,
            I => \N__28118\
        );

    \I__4789\ : Span4Mux_h
    port map (
            O => \N__28160\,
            I => \N__28115\
        );

    \I__4788\ : Span4Mux_h
    port map (
            O => \N__28157\,
            I => \N__28106\
        );

    \I__4787\ : Span4Mux_v
    port map (
            O => \N__28150\,
            I => \N__28106\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__28147\,
            I => \N__28106\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__28140\,
            I => \N__28106\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__28127\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__28118\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4782\ : Odrv4
    port map (
            O => \N__28115\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__28106\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4780\ : CascadeMux
    port map (
            O => \N__28097\,
            I => \N__28094\
        );

    \I__4779\ : InMux
    port map (
            O => \N__28094\,
            I => \N__28091\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__28091\,
            I => \N__28087\
        );

    \I__4777\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28083\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__28087\,
            I => \N__28080\
        );

    \I__4775\ : InMux
    port map (
            O => \N__28086\,
            I => \N__28077\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__28083\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__28080\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__28077\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__28070\,
            I => \N__28057\
        );

    \I__4770\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28049\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28068\,
            I => \N__28049\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28067\,
            I => \N__28049\
        );

    \I__4767\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28046\
        );

    \I__4766\ : InMux
    port map (
            O => \N__28065\,
            I => \N__28039\
        );

    \I__4765\ : InMux
    port map (
            O => \N__28064\,
            I => \N__28039\
        );

    \I__4764\ : InMux
    port map (
            O => \N__28063\,
            I => \N__28039\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28062\,
            I => \N__28028\
        );

    \I__4762\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28028\
        );

    \I__4761\ : InMux
    port map (
            O => \N__28060\,
            I => \N__28028\
        );

    \I__4760\ : InMux
    port map (
            O => \N__28057\,
            I => \N__28028\
        );

    \I__4759\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28028\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__28049\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__28046\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__28039\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__28028\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__4754\ : InMux
    port map (
            O => \N__28019\,
            I => \N__28015\
        );

    \I__4753\ : InMux
    port map (
            O => \N__28018\,
            I => \N__28012\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28015\,
            I => \elapsed_time_ns_1_RNIP3OD11_0_30\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__28012\,
            I => \elapsed_time_ns_1_RNIP3OD11_0_30\
        );

    \I__4750\ : InMux
    port map (
            O => \N__28007\,
            I => \N__28003\
        );

    \I__4749\ : InMux
    port map (
            O => \N__28006\,
            I => \N__28000\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__28003\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__28000\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__27995\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31_cascade_\
        );

    \I__4745\ : InMux
    port map (
            O => \N__27992\,
            I => \N__27988\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__27991\,
            I => \N__27985\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__27988\,
            I => \N__27981\
        );

    \I__4742\ : InMux
    port map (
            O => \N__27985\,
            I => \N__27978\
        );

    \I__4741\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27975\
        );

    \I__4740\ : Span4Mux_h
    port map (
            O => \N__27981\,
            I => \N__27972\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__27978\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__27975\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\
        );

    \I__4737\ : Odrv4
    port map (
            O => \N__27972\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__27965\,
            I => \N__27961\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__27964\,
            I => \N__27954\
        );

    \I__4734\ : InMux
    port map (
            O => \N__27961\,
            I => \N__27947\
        );

    \I__4733\ : InMux
    port map (
            O => \N__27960\,
            I => \N__27947\
        );

    \I__4732\ : InMux
    port map (
            O => \N__27959\,
            I => \N__27947\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__27958\,
            I => \N__27943\
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__27957\,
            I => \N__27940\
        );

    \I__4729\ : InMux
    port map (
            O => \N__27954\,
            I => \N__27936\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__27947\,
            I => \N__27933\
        );

    \I__4727\ : InMux
    port map (
            O => \N__27946\,
            I => \N__27928\
        );

    \I__4726\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27928\
        );

    \I__4725\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27925\
        );

    \I__4724\ : InMux
    port map (
            O => \N__27939\,
            I => \N__27922\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__27936\,
            I => \N__27917\
        );

    \I__4722\ : Span4Mux_h
    port map (
            O => \N__27933\,
            I => \N__27917\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__27928\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__27925\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__27922\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10\
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__27917\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10\
        );

    \I__4717\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27904\
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__27907\,
            I => \N__27901\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__27904\,
            I => \N__27898\
        );

    \I__4714\ : InMux
    port map (
            O => \N__27901\,
            I => \N__27893\
        );

    \I__4713\ : Span4Mux_v
    port map (
            O => \N__27898\,
            I => \N__27890\
        );

    \I__4712\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27885\
        );

    \I__4711\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27885\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__27893\,
            I => \elapsed_time_ns_1_RNIQ2MD11_0_13\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__27890\,
            I => \elapsed_time_ns_1_RNIQ2MD11_0_13\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__27885\,
            I => \elapsed_time_ns_1_RNIQ2MD11_0_13\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__27878\,
            I => \N__27875\
        );

    \I__4706\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27858\
        );

    \I__4705\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27841\
        );

    \I__4704\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27841\
        );

    \I__4703\ : InMux
    port map (
            O => \N__27872\,
            I => \N__27841\
        );

    \I__4702\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27841\
        );

    \I__4701\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27830\
        );

    \I__4700\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27830\
        );

    \I__4699\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27830\
        );

    \I__4698\ : InMux
    port map (
            O => \N__27867\,
            I => \N__27830\
        );

    \I__4697\ : InMux
    port map (
            O => \N__27866\,
            I => \N__27830\
        );

    \I__4696\ : InMux
    port map (
            O => \N__27865\,
            I => \N__27819\
        );

    \I__4695\ : InMux
    port map (
            O => \N__27864\,
            I => \N__27819\
        );

    \I__4694\ : InMux
    port map (
            O => \N__27863\,
            I => \N__27819\
        );

    \I__4693\ : InMux
    port map (
            O => \N__27862\,
            I => \N__27819\
        );

    \I__4692\ : InMux
    port map (
            O => \N__27861\,
            I => \N__27819\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__27858\,
            I => \N__27816\
        );

    \I__4690\ : CascadeMux
    port map (
            O => \N__27857\,
            I => \N__27812\
        );

    \I__4689\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27807\
        );

    \I__4688\ : InMux
    port map (
            O => \N__27855\,
            I => \N__27794\
        );

    \I__4687\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27794\
        );

    \I__4686\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27794\
        );

    \I__4685\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27794\
        );

    \I__4684\ : InMux
    port map (
            O => \N__27851\,
            I => \N__27794\
        );

    \I__4683\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27794\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__27841\,
            I => \N__27791\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__27830\,
            I => \N__27784\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__27819\,
            I => \N__27784\
        );

    \I__4679\ : Span4Mux_h
    port map (
            O => \N__27816\,
            I => \N__27784\
        );

    \I__4678\ : InMux
    port map (
            O => \N__27815\,
            I => \N__27777\
        );

    \I__4677\ : InMux
    port map (
            O => \N__27812\,
            I => \N__27777\
        );

    \I__4676\ : InMux
    port map (
            O => \N__27811\,
            I => \N__27777\
        );

    \I__4675\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27774\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__27807\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__27794\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__27791\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4671\ : Odrv4
    port map (
            O => \N__27784\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__27777\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__27774\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__27761\,
            I => \N__27757\
        );

    \I__4667\ : InMux
    port map (
            O => \N__27760\,
            I => \N__27754\
        );

    \I__4666\ : InMux
    port map (
            O => \N__27757\,
            I => \N__27748\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__27754\,
            I => \N__27745\
        );

    \I__4664\ : InMux
    port map (
            O => \N__27753\,
            I => \N__27741\
        );

    \I__4663\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27738\
        );

    \I__4662\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27735\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__27748\,
            I => \N__27732\
        );

    \I__4660\ : Span4Mux_h
    port map (
            O => \N__27745\,
            I => \N__27729\
        );

    \I__4659\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27726\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__27741\,
            I => \N__27723\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__27738\,
            I => \N__27718\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27718\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__27732\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__4654\ : Odrv4
    port map (
            O => \N__27729\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__27726\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__27723\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__4651\ : Odrv4
    port map (
            O => \N__27718\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__4650\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27703\
        );

    \I__4649\ : InMux
    port map (
            O => \N__27706\,
            I => \N__27698\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__27703\,
            I => \N__27695\
        );

    \I__4647\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27692\
        );

    \I__4646\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27689\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__27698\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7\
        );

    \I__4644\ : Odrv4
    port map (
            O => \N__27695\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__27692\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__27689\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7\
        );

    \I__4641\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27674\
        );

    \I__4640\ : CascadeMux
    port map (
            O => \N__27679\,
            I => \N__27671\
        );

    \I__4639\ : InMux
    port map (
            O => \N__27678\,
            I => \N__27668\
        );

    \I__4638\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27665\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__27674\,
            I => \N__27662\
        );

    \I__4636\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27659\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__27668\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__27665\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4633\ : Odrv4
    port map (
            O => \N__27662\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__27659\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4631\ : CascadeMux
    port map (
            O => \N__27650\,
            I => \N__27646\
        );

    \I__4630\ : CascadeMux
    port map (
            O => \N__27649\,
            I => \N__27643\
        );

    \I__4629\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27640\
        );

    \I__4628\ : InMux
    port map (
            O => \N__27643\,
            I => \N__27637\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__27640\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__27637\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\
        );

    \I__4625\ : CascadeMux
    port map (
            O => \N__27632\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\
        );

    \I__4624\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27623\
        );

    \I__4623\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27623\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__27623\,
            I => \N__27619\
        );

    \I__4621\ : InMux
    port map (
            O => \N__27622\,
            I => \N__27616\
        );

    \I__4620\ : Odrv12
    port map (
            O => \N__27619\,
            I => \elapsed_time_ns_1_RNIDP2KD1_0_1\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__27616\,
            I => \elapsed_time_ns_1_RNIDP2KD1_0_1\
        );

    \I__4618\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27608\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__27608\,
            I => \N__27605\
        );

    \I__4616\ : Odrv4
    port map (
            O => \N__27605\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\
        );

    \I__4615\ : CascadeMux
    port map (
            O => \N__27602\,
            I => \elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_\
        );

    \I__4614\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27595\
        );

    \I__4613\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27592\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__27595\,
            I => \phase_controller_inst1.stoper_hc.N_307\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__27592\,
            I => \phase_controller_inst1.stoper_hc.N_307\
        );

    \I__4610\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27583\
        );

    \I__4609\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27580\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__27583\,
            I => \N__27576\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__27580\,
            I => \N__27573\
        );

    \I__4606\ : InMux
    port map (
            O => \N__27579\,
            I => \N__27570\
        );

    \I__4605\ : Odrv12
    port map (
            O => \N__27576\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__4604\ : Odrv12
    port map (
            O => \N__27573\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__27570\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__4602\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27560\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__27560\,
            I => \N__27557\
        );

    \I__4600\ : Odrv4
    port map (
            O => \N__27557\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_10\
        );

    \I__4599\ : CascadeMux
    port map (
            O => \N__27554\,
            I => \N__27551\
        );

    \I__4598\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27548\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__27548\,
            I => \N__27545\
        );

    \I__4596\ : Span4Mux_h
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__27542\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\
        );

    \I__4594\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27536\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__27536\,
            I => \N__27533\
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__27533\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__27530\,
            I => \N__27525\
        );

    \I__4590\ : CascadeMux
    port map (
            O => \N__27529\,
            I => \N__27522\
        );

    \I__4589\ : CascadeMux
    port map (
            O => \N__27528\,
            I => \N__27519\
        );

    \I__4588\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27516\
        );

    \I__4587\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27511\
        );

    \I__4586\ : InMux
    port map (
            O => \N__27519\,
            I => \N__27511\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__27516\,
            I => \N__27506\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__27511\,
            I => \N__27503\
        );

    \I__4583\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27500\
        );

    \I__4582\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27497\
        );

    \I__4581\ : Span12Mux_v
    port map (
            O => \N__27506\,
            I => \N__27494\
        );

    \I__4580\ : Span4Mux_h
    port map (
            O => \N__27503\,
            I => \N__27491\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__27500\,
            I => \N__27488\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__27497\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4577\ : Odrv12
    port map (
            O => \N__27494\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__27491\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4575\ : Odrv12
    port map (
            O => \N__27488\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4574\ : CascadeMux
    port map (
            O => \N__27479\,
            I => \N__27476\
        );

    \I__4573\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27473\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__27473\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__4571\ : InMux
    port map (
            O => \N__27470\,
            I => \N__27467\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__27467\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__4569\ : InMux
    port map (
            O => \N__27464\,
            I => \N__27461\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__27461\,
            I => \N__27455\
        );

    \I__4567\ : InMux
    port map (
            O => \N__27460\,
            I => \N__27452\
        );

    \I__4566\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27449\
        );

    \I__4565\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27446\
        );

    \I__4564\ : Span4Mux_v
    port map (
            O => \N__27455\,
            I => \N__27443\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__27452\,
            I => \N__27440\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__27449\,
            I => \N__27435\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__27446\,
            I => \N__27435\
        );

    \I__4560\ : Span4Mux_h
    port map (
            O => \N__27443\,
            I => \N__27432\
        );

    \I__4559\ : Span4Mux_h
    port map (
            O => \N__27440\,
            I => \N__27429\
        );

    \I__4558\ : Span4Mux_h
    port map (
            O => \N__27435\,
            I => \N__27426\
        );

    \I__4557\ : Odrv4
    port map (
            O => \N__27432\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4556\ : Odrv4
    port map (
            O => \N__27429\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4555\ : Odrv4
    port map (
            O => \N__27426\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__27419\,
            I => \N__27416\
        );

    \I__4553\ : InMux
    port map (
            O => \N__27416\,
            I => \N__27413\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__27413\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__4551\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27407\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__27407\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27392\
        );

    \I__4548\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27380\
        );

    \I__4547\ : InMux
    port map (
            O => \N__27402\,
            I => \N__27380\
        );

    \I__4546\ : InMux
    port map (
            O => \N__27401\,
            I => \N__27380\
        );

    \I__4545\ : InMux
    port map (
            O => \N__27400\,
            I => \N__27359\
        );

    \I__4544\ : InMux
    port map (
            O => \N__27399\,
            I => \N__27359\
        );

    \I__4543\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27359\
        );

    \I__4542\ : InMux
    port map (
            O => \N__27397\,
            I => \N__27359\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27396\,
            I => \N__27359\
        );

    \I__4540\ : InMux
    port map (
            O => \N__27395\,
            I => \N__27356\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__27392\,
            I => \N__27353\
        );

    \I__4538\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27342\
        );

    \I__4537\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27342\
        );

    \I__4536\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27342\
        );

    \I__4535\ : InMux
    port map (
            O => \N__27388\,
            I => \N__27342\
        );

    \I__4534\ : InMux
    port map (
            O => \N__27387\,
            I => \N__27342\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__27380\,
            I => \N__27339\
        );

    \I__4532\ : InMux
    port map (
            O => \N__27379\,
            I => \N__27328\
        );

    \I__4531\ : InMux
    port map (
            O => \N__27378\,
            I => \N__27328\
        );

    \I__4530\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27328\
        );

    \I__4529\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27328\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27375\,
            I => \N__27328\
        );

    \I__4527\ : InMux
    port map (
            O => \N__27374\,
            I => \N__27311\
        );

    \I__4526\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27311\
        );

    \I__4525\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27311\
        );

    \I__4524\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27311\
        );

    \I__4523\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27311\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__27359\,
            I => \N__27305\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__27356\,
            I => \N__27305\
        );

    \I__4520\ : Span4Mux_v
    port map (
            O => \N__27353\,
            I => \N__27302\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__27342\,
            I => \N__27295\
        );

    \I__4518\ : Span4Mux_h
    port map (
            O => \N__27339\,
            I => \N__27295\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__27328\,
            I => \N__27295\
        );

    \I__4516\ : InMux
    port map (
            O => \N__27327\,
            I => \N__27282\
        );

    \I__4515\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27282\
        );

    \I__4514\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27282\
        );

    \I__4513\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27282\
        );

    \I__4512\ : InMux
    port map (
            O => \N__27323\,
            I => \N__27282\
        );

    \I__4511\ : InMux
    port map (
            O => \N__27322\,
            I => \N__27282\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__27311\,
            I => \N__27279\
        );

    \I__4509\ : InMux
    port map (
            O => \N__27310\,
            I => \N__27276\
        );

    \I__4508\ : Span4Mux_v
    port map (
            O => \N__27305\,
            I => \N__27273\
        );

    \I__4507\ : Span4Mux_h
    port map (
            O => \N__27302\,
            I => \N__27268\
        );

    \I__4506\ : Span4Mux_v
    port map (
            O => \N__27295\,
            I => \N__27268\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__27282\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4504\ : Odrv4
    port map (
            O => \N__27279\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__27276\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4502\ : Odrv4
    port map (
            O => \N__27273\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4501\ : Odrv4
    port map (
            O => \N__27268\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4500\ : CascadeMux
    port map (
            O => \N__27257\,
            I => \N__27244\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__27256\,
            I => \N__27241\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27255\,
            I => \N__27225\
        );

    \I__4497\ : InMux
    port map (
            O => \N__27254\,
            I => \N__27225\
        );

    \I__4496\ : InMux
    port map (
            O => \N__27253\,
            I => \N__27225\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27225\
        );

    \I__4494\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27225\
        );

    \I__4493\ : InMux
    port map (
            O => \N__27250\,
            I => \N__27225\
        );

    \I__4492\ : InMux
    port map (
            O => \N__27249\,
            I => \N__27210\
        );

    \I__4491\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27210\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27247\,
            I => \N__27210\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27210\
        );

    \I__4488\ : InMux
    port map (
            O => \N__27241\,
            I => \N__27210\
        );

    \I__4487\ : InMux
    port map (
            O => \N__27240\,
            I => \N__27203\
        );

    \I__4486\ : InMux
    port map (
            O => \N__27239\,
            I => \N__27203\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27238\,
            I => \N__27203\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27225\,
            I => \N__27190\
        );

    \I__4483\ : InMux
    port map (
            O => \N__27224\,
            I => \N__27181\
        );

    \I__4482\ : InMux
    port map (
            O => \N__27223\,
            I => \N__27181\
        );

    \I__4481\ : InMux
    port map (
            O => \N__27222\,
            I => \N__27181\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27221\,
            I => \N__27181\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__27210\,
            I => \N__27178\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__27203\,
            I => \N__27175\
        );

    \I__4477\ : InMux
    port map (
            O => \N__27202\,
            I => \N__27164\
        );

    \I__4476\ : InMux
    port map (
            O => \N__27201\,
            I => \N__27164\
        );

    \I__4475\ : InMux
    port map (
            O => \N__27200\,
            I => \N__27164\
        );

    \I__4474\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27164\
        );

    \I__4473\ : InMux
    port map (
            O => \N__27198\,
            I => \N__27164\
        );

    \I__4472\ : InMux
    port map (
            O => \N__27197\,
            I => \N__27153\
        );

    \I__4471\ : InMux
    port map (
            O => \N__27196\,
            I => \N__27153\
        );

    \I__4470\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27153\
        );

    \I__4469\ : InMux
    port map (
            O => \N__27194\,
            I => \N__27153\
        );

    \I__4468\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27153\
        );

    \I__4467\ : Span4Mux_v
    port map (
            O => \N__27190\,
            I => \N__27150\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__27181\,
            I => \N__27143\
        );

    \I__4465\ : Span4Mux_h
    port map (
            O => \N__27178\,
            I => \N__27143\
        );

    \I__4464\ : Span4Mux_v
    port map (
            O => \N__27175\,
            I => \N__27143\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__27164\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27153\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__27150\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4460\ : Odrv4
    port map (
            O => \N__27143\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__27134\,
            I => \N__27131\
        );

    \I__4458\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27128\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__27128\,
            I => \N__27125\
        );

    \I__4456\ : Span4Mux_v
    port map (
            O => \N__27125\,
            I => \N__27122\
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__27122\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__4454\ : CascadeMux
    port map (
            O => \N__27119\,
            I => \N__27106\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__27118\,
            I => \N__27103\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__27117\,
            I => \N__27100\
        );

    \I__4451\ : CascadeMux
    port map (
            O => \N__27116\,
            I => \N__27095\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__27115\,
            I => \N__27085\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__27114\,
            I => \N__27077\
        );

    \I__4448\ : CascadeMux
    port map (
            O => \N__27113\,
            I => \N__27074\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__27112\,
            I => \N__27071\
        );

    \I__4446\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27056\
        );

    \I__4445\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27056\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27109\,
            I => \N__27056\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27106\,
            I => \N__27056\
        );

    \I__4442\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27056\
        );

    \I__4441\ : InMux
    port map (
            O => \N__27100\,
            I => \N__27056\
        );

    \I__4440\ : InMux
    port map (
            O => \N__27099\,
            I => \N__27049\
        );

    \I__4439\ : InMux
    port map (
            O => \N__27098\,
            I => \N__27049\
        );

    \I__4438\ : InMux
    port map (
            O => \N__27095\,
            I => \N__27049\
        );

    \I__4437\ : CascadeMux
    port map (
            O => \N__27094\,
            I => \N__27044\
        );

    \I__4436\ : CascadeMux
    port map (
            O => \N__27093\,
            I => \N__27041\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__27092\,
            I => \N__27038\
        );

    \I__4434\ : CascadeMux
    port map (
            O => \N__27091\,
            I => \N__27032\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__27090\,
            I => \N__27029\
        );

    \I__4432\ : InMux
    port map (
            O => \N__27089\,
            I => \N__27024\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27024\
        );

    \I__4430\ : InMux
    port map (
            O => \N__27085\,
            I => \N__27021\
        );

    \I__4429\ : InMux
    port map (
            O => \N__27084\,
            I => \N__27010\
        );

    \I__4428\ : InMux
    port map (
            O => \N__27083\,
            I => \N__27010\
        );

    \I__4427\ : InMux
    port map (
            O => \N__27082\,
            I => \N__27010\
        );

    \I__4426\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27010\
        );

    \I__4425\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27010\
        );

    \I__4424\ : InMux
    port map (
            O => \N__27077\,
            I => \N__27003\
        );

    \I__4423\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27003\
        );

    \I__4422\ : InMux
    port map (
            O => \N__27071\,
            I => \N__27003\
        );

    \I__4421\ : InMux
    port map (
            O => \N__27070\,
            I => \N__26998\
        );

    \I__4420\ : InMux
    port map (
            O => \N__27069\,
            I => \N__26998\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__27056\,
            I => \N__26995\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__27049\,
            I => \N__26992\
        );

    \I__4417\ : InMux
    port map (
            O => \N__27048\,
            I => \N__26981\
        );

    \I__4416\ : InMux
    port map (
            O => \N__27047\,
            I => \N__26981\
        );

    \I__4415\ : InMux
    port map (
            O => \N__27044\,
            I => \N__26981\
        );

    \I__4414\ : InMux
    port map (
            O => \N__27041\,
            I => \N__26981\
        );

    \I__4413\ : InMux
    port map (
            O => \N__27038\,
            I => \N__26981\
        );

    \I__4412\ : InMux
    port map (
            O => \N__27037\,
            I => \N__26970\
        );

    \I__4411\ : InMux
    port map (
            O => \N__27036\,
            I => \N__26970\
        );

    \I__4410\ : InMux
    port map (
            O => \N__27035\,
            I => \N__26970\
        );

    \I__4409\ : InMux
    port map (
            O => \N__27032\,
            I => \N__26970\
        );

    \I__4408\ : InMux
    port map (
            O => \N__27029\,
            I => \N__26970\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__26959\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__27021\,
            I => \N__26959\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__27010\,
            I => \N__26959\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__27003\,
            I => \N__26959\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__26998\,
            I => \N__26959\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__26995\,
            I => \N__26956\
        );

    \I__4401\ : Span4Mux_h
    port map (
            O => \N__26992\,
            I => \N__26953\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__26981\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__26970\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__4398\ : Odrv12
    port map (
            O => \N__26959\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__26956\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__4396\ : Odrv4
    port map (
            O => \N__26953\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__4395\ : CascadeMux
    port map (
            O => \N__26942\,
            I => \N__26939\
        );

    \I__4394\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26934\
        );

    \I__4393\ : CascadeMux
    port map (
            O => \N__26938\,
            I => \N__26931\
        );

    \I__4392\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26927\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__26934\,
            I => \N__26924\
        );

    \I__4390\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26921\
        );

    \I__4389\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26918\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__26927\,
            I => \N__26915\
        );

    \I__4387\ : Span4Mux_v
    port map (
            O => \N__26924\,
            I => \N__26910\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__26921\,
            I => \N__26910\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__26918\,
            I => \N__26903\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__26915\,
            I => \N__26903\
        );

    \I__4383\ : Span4Mux_h
    port map (
            O => \N__26910\,
            I => \N__26903\
        );

    \I__4382\ : Span4Mux_v
    port map (
            O => \N__26903\,
            I => \N__26899\
        );

    \I__4381\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26896\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__26899\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__26896\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__26891\,
            I => \N__26887\
        );

    \I__4377\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26884\
        );

    \I__4376\ : InMux
    port map (
            O => \N__26887\,
            I => \N__26879\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__26884\,
            I => \N__26876\
        );

    \I__4374\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26871\
        );

    \I__4373\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26871\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__26879\,
            I => \elapsed_time_ns_1_RNIO0MD11_0_11\
        );

    \I__4371\ : Odrv4
    port map (
            O => \N__26876\,
            I => \elapsed_time_ns_1_RNIO0MD11_0_11\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__26871\,
            I => \elapsed_time_ns_1_RNIO0MD11_0_11\
        );

    \I__4369\ : CascadeMux
    port map (
            O => \N__26864\,
            I => \N__26860\
        );

    \I__4368\ : InMux
    port map (
            O => \N__26863\,
            I => \N__26857\
        );

    \I__4367\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26854\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__26857\,
            I => \N__26851\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__26854\,
            I => \N__26848\
        );

    \I__4364\ : Span4Mux_h
    port map (
            O => \N__26851\,
            I => \N__26842\
        );

    \I__4363\ : Span4Mux_v
    port map (
            O => \N__26848\,
            I => \N__26842\
        );

    \I__4362\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26839\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__26842\,
            I => \elapsed_time_ns_1_RNIP1MD11_0_12\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__26839\,
            I => \elapsed_time_ns_1_RNIP1MD11_0_12\
        );

    \I__4359\ : InMux
    port map (
            O => \N__26834\,
            I => \N__26831\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__26831\,
            I => \current_shift_inst.PI_CTRL.integrator_i_10\
        );

    \I__4357\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26825\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__26825\,
            I => \N__26822\
        );

    \I__4355\ : Odrv12
    port map (
            O => \N__26822\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__26819\,
            I => \N__26816\
        );

    \I__4353\ : InMux
    port map (
            O => \N__26816\,
            I => \N__26812\
        );

    \I__4352\ : InMux
    port map (
            O => \N__26815\,
            I => \N__26808\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__26812\,
            I => \N__26805\
        );

    \I__4350\ : InMux
    port map (
            O => \N__26811\,
            I => \N__26800\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__26808\,
            I => \N__26797\
        );

    \I__4348\ : Span4Mux_h
    port map (
            O => \N__26805\,
            I => \N__26794\
        );

    \I__4347\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26791\
        );

    \I__4346\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26788\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__26800\,
            I => \N__26785\
        );

    \I__4344\ : Span4Mux_h
    port map (
            O => \N__26797\,
            I => \N__26778\
        );

    \I__4343\ : Span4Mux_h
    port map (
            O => \N__26794\,
            I => \N__26778\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__26791\,
            I => \N__26778\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__26788\,
            I => \N__26775\
        );

    \I__4340\ : Odrv12
    port map (
            O => \N__26785\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__26778\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__26775\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4337\ : InMux
    port map (
            O => \N__26768\,
            I => \N__26765\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__26765\,
            I => \N__26762\
        );

    \I__4335\ : Odrv4
    port map (
            O => \N__26762\,
            I => \current_shift_inst.PI_CTRL.integrator_i_20\
        );

    \I__4334\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26755\
        );

    \I__4333\ : InMux
    port map (
            O => \N__26758\,
            I => \N__26751\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__26755\,
            I => \N__26748\
        );

    \I__4331\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26745\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__26751\,
            I => \N__26742\
        );

    \I__4329\ : Span4Mux_h
    port map (
            O => \N__26748\,
            I => \N__26739\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__26745\,
            I => \N__26736\
        );

    \I__4327\ : Odrv12
    port map (
            O => \N__26742\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__26739\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__4325\ : Odrv12
    port map (
            O => \N__26736\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__4324\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26726\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__26726\,
            I => \N__26723\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__26723\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\
        );

    \I__4321\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26717\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__26717\,
            I => \N__26714\
        );

    \I__4319\ : Odrv12
    port map (
            O => \N__26714\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__4318\ : InMux
    port map (
            O => \N__26711\,
            I => \N__26707\
        );

    \I__4317\ : InMux
    port map (
            O => \N__26710\,
            I => \N__26704\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__26707\,
            I => \N__26698\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__26704\,
            I => \N__26698\
        );

    \I__4314\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26695\
        );

    \I__4313\ : Span4Mux_v
    port map (
            O => \N__26698\,
            I => \N__26692\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__26695\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__4311\ : Odrv4
    port map (
            O => \N__26692\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__26687\,
            I => \N__26684\
        );

    \I__4309\ : InMux
    port map (
            O => \N__26684\,
            I => \N__26681\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__26681\,
            I => \N__26675\
        );

    \I__4307\ : InMux
    port map (
            O => \N__26680\,
            I => \N__26672\
        );

    \I__4306\ : InMux
    port map (
            O => \N__26679\,
            I => \N__26669\
        );

    \I__4305\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26665\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__26675\,
            I => \N__26658\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__26672\,
            I => \N__26658\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__26669\,
            I => \N__26658\
        );

    \I__4301\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26655\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__26665\,
            I => \N__26650\
        );

    \I__4299\ : Span4Mux_h
    port map (
            O => \N__26658\,
            I => \N__26650\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__26655\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__4297\ : Odrv4
    port map (
            O => \N__26650\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__4296\ : InMux
    port map (
            O => \N__26645\,
            I => \N__26642\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__26642\,
            I => \N__26639\
        );

    \I__4294\ : Span4Mux_v
    port map (
            O => \N__26639\,
            I => \N__26634\
        );

    \I__4293\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26631\
        );

    \I__4292\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26628\
        );

    \I__4291\ : Span4Mux_h
    port map (
            O => \N__26634\,
            I => \N__26625\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__26631\,
            I => \N__26622\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__26628\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__4288\ : Odrv4
    port map (
            O => \N__26625\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__4287\ : Odrv12
    port map (
            O => \N__26622\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__4286\ : InMux
    port map (
            O => \N__26615\,
            I => \N__26612\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__26612\,
            I => \N__26609\
        );

    \I__4284\ : Span4Mux_h
    port map (
            O => \N__26609\,
            I => \N__26606\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__26606\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__26603\,
            I => \N__26600\
        );

    \I__4281\ : InMux
    port map (
            O => \N__26600\,
            I => \N__26597\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__26597\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\
        );

    \I__4279\ : InMux
    port map (
            O => \N__26594\,
            I => \N__26590\
        );

    \I__4278\ : InMux
    port map (
            O => \N__26593\,
            I => \N__26587\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__26590\,
            I => \N__26583\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__26587\,
            I => \N__26580\
        );

    \I__4275\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26577\
        );

    \I__4274\ : Span4Mux_h
    port map (
            O => \N__26583\,
            I => \N__26574\
        );

    \I__4273\ : Span4Mux_v
    port map (
            O => \N__26580\,
            I => \N__26571\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__26577\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__26574\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__26571\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__4269\ : CascadeMux
    port map (
            O => \N__26564\,
            I => \N__26560\
        );

    \I__4268\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26556\
        );

    \I__4267\ : InMux
    port map (
            O => \N__26560\,
            I => \N__26553\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__26559\,
            I => \N__26550\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__26556\,
            I => \N__26546\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__26553\,
            I => \N__26543\
        );

    \I__4263\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26540\
        );

    \I__4262\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26537\
        );

    \I__4261\ : Span4Mux_h
    port map (
            O => \N__26546\,
            I => \N__26534\
        );

    \I__4260\ : Span4Mux_v
    port map (
            O => \N__26543\,
            I => \N__26528\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__26540\,
            I => \N__26528\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__26537\,
            I => \N__26523\
        );

    \I__4257\ : Span4Mux_h
    port map (
            O => \N__26534\,
            I => \N__26523\
        );

    \I__4256\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26520\
        );

    \I__4255\ : Span4Mux_h
    port map (
            O => \N__26528\,
            I => \N__26517\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__26523\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__26520\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4252\ : Odrv4
    port map (
            O => \N__26517\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__26510\,
            I => \N__26507\
        );

    \I__4250\ : InMux
    port map (
            O => \N__26507\,
            I => \N__26504\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__26504\,
            I => \N__26501\
        );

    \I__4248\ : Span4Mux_h
    port map (
            O => \N__26501\,
            I => \N__26498\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__26498\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\
        );

    \I__4246\ : CascadeMux
    port map (
            O => \N__26495\,
            I => \N__26492\
        );

    \I__4245\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26489\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__26489\,
            I => \N__26486\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__26486\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\
        );

    \I__4242\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26480\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__26480\,
            I => \N__26477\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__26477\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__26474\,
            I => \N__26471\
        );

    \I__4238\ : InMux
    port map (
            O => \N__26471\,
            I => \N__26468\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__26468\,
            I => \N__26465\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__26465\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__4235\ : InMux
    port map (
            O => \N__26462\,
            I => \N__26457\
        );

    \I__4234\ : InMux
    port map (
            O => \N__26461\,
            I => \N__26454\
        );

    \I__4233\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26451\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__26457\,
            I => \N__26448\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__26454\,
            I => \N__26445\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__26451\,
            I => \N__26442\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__26448\,
            I => \N__26439\
        );

    \I__4228\ : Span4Mux_h
    port map (
            O => \N__26445\,
            I => \N__26436\
        );

    \I__4227\ : Span4Mux_h
    port map (
            O => \N__26442\,
            I => \N__26433\
        );

    \I__4226\ : Odrv4
    port map (
            O => \N__26439\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__26436\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__4224\ : Odrv4
    port map (
            O => \N__26433\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__4223\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26423\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__4221\ : Span4Mux_h
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__26417\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__26414\,
            I => \N__26411\
        );

    \I__4218\ : InMux
    port map (
            O => \N__26411\,
            I => \N__26407\
        );

    \I__4217\ : InMux
    port map (
            O => \N__26410\,
            I => \N__26404\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__26407\,
            I => \N__26401\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__26404\,
            I => \N__26397\
        );

    \I__4214\ : Span4Mux_h
    port map (
            O => \N__26401\,
            I => \N__26394\
        );

    \I__4213\ : InMux
    port map (
            O => \N__26400\,
            I => \N__26390\
        );

    \I__4212\ : Span4Mux_h
    port map (
            O => \N__26397\,
            I => \N__26387\
        );

    \I__4211\ : Span4Mux_h
    port map (
            O => \N__26394\,
            I => \N__26384\
        );

    \I__4210\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26381\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__26390\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4208\ : Odrv4
    port map (
            O => \N__26387\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4207\ : Odrv4
    port map (
            O => \N__26384\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__26381\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__26372\,
            I => \N__26369\
        );

    \I__4204\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__26366\,
            I => \current_shift_inst.PI_CTRL.integrator_i_1\
        );

    \I__4202\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26360\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__26360\,
            I => \current_shift_inst.PI_CTRL.integrator_i_21\
        );

    \I__4200\ : CascadeMux
    port map (
            O => \N__26357\,
            I => \N__26354\
        );

    \I__4199\ : InMux
    port map (
            O => \N__26354\,
            I => \N__26350\
        );

    \I__4198\ : InMux
    port map (
            O => \N__26353\,
            I => \N__26347\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__26350\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_12\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__26347\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_12\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__26342\,
            I => \N__26339\
        );

    \I__4194\ : InMux
    port map (
            O => \N__26339\,
            I => \N__26335\
        );

    \I__4193\ : InMux
    port map (
            O => \N__26338\,
            I => \N__26332\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__26335\,
            I => \N__26328\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__26332\,
            I => \N__26323\
        );

    \I__4190\ : InMux
    port map (
            O => \N__26331\,
            I => \N__26320\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__26328\,
            I => \N__26317\
        );

    \I__4188\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26312\
        );

    \I__4187\ : InMux
    port map (
            O => \N__26326\,
            I => \N__26312\
        );

    \I__4186\ : Span4Mux_h
    port map (
            O => \N__26323\,
            I => \N__26309\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__26320\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__26317\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__26312\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__26309\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4181\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26297\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__26297\,
            I => \current_shift_inst.PI_CTRL.integrator_i_14\
        );

    \I__4179\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26291\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__26291\,
            I => \current_shift_inst.PI_CTRL.integrator_i_22\
        );

    \I__4177\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26284\
        );

    \I__4176\ : InMux
    port map (
            O => \N__26287\,
            I => \N__26280\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__26284\,
            I => \N__26277\
        );

    \I__4174\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26274\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__26280\,
            I => \N__26269\
        );

    \I__4172\ : Span4Mux_h
    port map (
            O => \N__26277\,
            I => \N__26264\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__26274\,
            I => \N__26264\
        );

    \I__4170\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26261\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26272\,
            I => \N__26258\
        );

    \I__4168\ : Span4Mux_h
    port map (
            O => \N__26269\,
            I => \N__26253\
        );

    \I__4167\ : Span4Mux_h
    port map (
            O => \N__26264\,
            I => \N__26253\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__26261\,
            I => \N__26250\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__26258\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__4164\ : Odrv4
    port map (
            O => \N__26253\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__4163\ : Odrv12
    port map (
            O => \N__26250\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__4162\ : InMux
    port map (
            O => \N__26243\,
            I => \N__26240\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__26240\,
            I => \current_shift_inst.PI_CTRL.integrator_i_19\
        );

    \I__4160\ : InMux
    port map (
            O => \N__26237\,
            I => \N__26234\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__26234\,
            I => \N__26231\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__26231\,
            I => \current_shift_inst.PI_CTRL.integrator_i_6\
        );

    \I__4157\ : InMux
    port map (
            O => \N__26228\,
            I => \N__26225\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__4155\ : Span4Mux_v
    port map (
            O => \N__26222\,
            I => \N__26219\
        );

    \I__4154\ : Odrv4
    port map (
            O => \N__26219\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__26216\,
            I => \N__26213\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26213\,
            I => \N__26209\
        );

    \I__4151\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26206\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__26209\,
            I => \N__26203\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__26206\,
            I => \N__26199\
        );

    \I__4148\ : Span4Mux_h
    port map (
            O => \N__26203\,
            I => \N__26196\
        );

    \I__4147\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26193\
        );

    \I__4146\ : Odrv12
    port map (
            O => \N__26199\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__4145\ : Odrv4
    port map (
            O => \N__26196\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__26193\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__4143\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26183\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26180\
        );

    \I__4141\ : Span4Mux_h
    port map (
            O => \N__26180\,
            I => \N__26177\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__26177\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_9\
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__26174\,
            I => \N__26171\
        );

    \I__4138\ : InMux
    port map (
            O => \N__26171\,
            I => \N__26168\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__26168\,
            I => \N__26165\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__26165\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\
        );

    \I__4135\ : CascadeMux
    port map (
            O => \N__26162\,
            I => \N__26159\
        );

    \I__4134\ : InMux
    port map (
            O => \N__26159\,
            I => \N__26156\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__26156\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__4132\ : CascadeMux
    port map (
            O => \N__26153\,
            I => \N__26150\
        );

    \I__4131\ : InMux
    port map (
            O => \N__26150\,
            I => \N__26146\
        );

    \I__4130\ : InMux
    port map (
            O => \N__26149\,
            I => \N__26143\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__26146\,
            I => \N__26139\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__26143\,
            I => \N__26135\
        );

    \I__4127\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26131\
        );

    \I__4126\ : Span4Mux_v
    port map (
            O => \N__26139\,
            I => \N__26128\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26125\
        );

    \I__4124\ : Span4Mux_h
    port map (
            O => \N__26135\,
            I => \N__26122\
        );

    \I__4123\ : InMux
    port map (
            O => \N__26134\,
            I => \N__26119\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__26131\,
            I => \N__26116\
        );

    \I__4121\ : Span4Mux_h
    port map (
            O => \N__26128\,
            I => \N__26111\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__26125\,
            I => \N__26111\
        );

    \I__4119\ : Span4Mux_h
    port map (
            O => \N__26122\,
            I => \N__26108\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__26119\,
            I => \N__26101\
        );

    \I__4117\ : Span4Mux_v
    port map (
            O => \N__26116\,
            I => \N__26101\
        );

    \I__4116\ : Span4Mux_h
    port map (
            O => \N__26111\,
            I => \N__26101\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__26108\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__26101\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4113\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26093\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26090\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__26090\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__26087\,
            I => \N__26084\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26084\,
            I => \N__26081\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__26081\,
            I => \N__26078\
        );

    \I__4107\ : Odrv4
    port map (
            O => \N__26078\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__4106\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26070\
        );

    \I__4105\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26067\
        );

    \I__4104\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26064\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__26070\,
            I => \N__26061\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__26067\,
            I => \N__26054\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__26064\,
            I => \N__26054\
        );

    \I__4100\ : Span4Mux_h
    port map (
            O => \N__26061\,
            I => \N__26054\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__26054\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__4098\ : InMux
    port map (
            O => \N__26051\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__4097\ : InMux
    port map (
            O => \N__26048\,
            I => \N__26044\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26047\,
            I => \N__26040\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__26044\,
            I => \N__26037\
        );

    \I__4094\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26034\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__26040\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__26037\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__26034\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26027\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__4089\ : InMux
    port map (
            O => \N__26024\,
            I => \N__26021\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__26021\,
            I => \N__26016\
        );

    \I__4087\ : InMux
    port map (
            O => \N__26020\,
            I => \N__26013\
        );

    \I__4086\ : InMux
    port map (
            O => \N__26019\,
            I => \N__26010\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__26016\,
            I => \N__26007\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__26013\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__26010\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__26007\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4081\ : InMux
    port map (
            O => \N__26000\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__4080\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25992\
        );

    \I__4079\ : InMux
    port map (
            O => \N__25996\,
            I => \N__25989\
        );

    \I__4078\ : InMux
    port map (
            O => \N__25995\,
            I => \N__25986\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__25992\,
            I => \N__25983\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__25989\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__25986\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4074\ : Odrv4
    port map (
            O => \N__25983\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4073\ : InMux
    port map (
            O => \N__25976\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__4072\ : InMux
    port map (
            O => \N__25973\,
            I => \N__25968\
        );

    \I__4071\ : InMux
    port map (
            O => \N__25972\,
            I => \N__25965\
        );

    \I__4070\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25962\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__25968\,
            I => \N__25959\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__25965\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__25962\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4066\ : Odrv12
    port map (
            O => \N__25959\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4065\ : InMux
    port map (
            O => \N__25952\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__4064\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25945\
        );

    \I__4063\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25941\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__25945\,
            I => \N__25938\
        );

    \I__4061\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25935\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__25941\,
            I => \N__25930\
        );

    \I__4059\ : Span4Mux_h
    port map (
            O => \N__25938\,
            I => \N__25930\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__25935\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4057\ : Odrv4
    port map (
            O => \N__25930\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4056\ : InMux
    port map (
            O => \N__25925\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__4055\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25917\
        );

    \I__4054\ : InMux
    port map (
            O => \N__25921\,
            I => \N__25914\
        );

    \I__4053\ : InMux
    port map (
            O => \N__25920\,
            I => \N__25911\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__25917\,
            I => \N__25908\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__25914\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__25911\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4049\ : Odrv4
    port map (
            O => \N__25908\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4048\ : InMux
    port map (
            O => \N__25901\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__4047\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25894\
        );

    \I__4046\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25890\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__25894\,
            I => \N__25887\
        );

    \I__4044\ : InMux
    port map (
            O => \N__25893\,
            I => \N__25884\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__25890\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__25887\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__25884\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4040\ : InMux
    port map (
            O => \N__25877\,
            I => \bfn_11_7_0_\
        );

    \I__4039\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25856\
        );

    \I__4038\ : InMux
    port map (
            O => \N__25873\,
            I => \N__25856\
        );

    \I__4037\ : InMux
    port map (
            O => \N__25872\,
            I => \N__25856\
        );

    \I__4036\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25856\
        );

    \I__4035\ : InMux
    port map (
            O => \N__25870\,
            I => \N__25851\
        );

    \I__4034\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25851\
        );

    \I__4033\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25842\
        );

    \I__4032\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25842\
        );

    \I__4031\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25842\
        );

    \I__4030\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25842\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__25856\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__25851\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__25842\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4026\ : InMux
    port map (
            O => \N__25835\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__4025\ : InMux
    port map (
            O => \N__25832\,
            I => \N__25828\
        );

    \I__4024\ : InMux
    port map (
            O => \N__25831\,
            I => \N__25824\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__25828\,
            I => \N__25821\
        );

    \I__4022\ : InMux
    port map (
            O => \N__25827\,
            I => \N__25818\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__25824\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4020\ : Odrv4
    port map (
            O => \N__25821\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__25818\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4018\ : InMux
    port map (
            O => \N__25811\,
            I => \N__25807\
        );

    \I__4017\ : InMux
    port map (
            O => \N__25810\,
            I => \N__25804\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__25807\,
            I => \N__25801\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__25804\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__25801\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4013\ : InMux
    port map (
            O => \N__25796\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__4012\ : InMux
    port map (
            O => \N__25793\,
            I => \N__25789\
        );

    \I__4011\ : InMux
    port map (
            O => \N__25792\,
            I => \N__25786\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__25789\,
            I => \N__25783\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__25786\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4008\ : Odrv4
    port map (
            O => \N__25783\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4007\ : InMux
    port map (
            O => \N__25778\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__4006\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25772\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__25772\,
            I => \N__25768\
        );

    \I__4004\ : InMux
    port map (
            O => \N__25771\,
            I => \N__25765\
        );

    \I__4003\ : Span4Mux_h
    port map (
            O => \N__25768\,
            I => \N__25762\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__25765\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4001\ : Odrv4
    port map (
            O => \N__25762\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4000\ : InMux
    port map (
            O => \N__25757\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__3999\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25750\
        );

    \I__3998\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25747\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__25750\,
            I => \N__25744\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__25747\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3995\ : Odrv12
    port map (
            O => \N__25744\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3994\ : InMux
    port map (
            O => \N__25739\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__3993\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25732\
        );

    \I__3992\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25729\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__25732\,
            I => \N__25726\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__25729\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__25726\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3988\ : InMux
    port map (
            O => \N__25721\,
            I => \bfn_10_26_0_\
        );

    \I__3987\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25714\
        );

    \I__3986\ : InMux
    port map (
            O => \N__25717\,
            I => \N__25711\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__25714\,
            I => \N__25708\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__25711\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3983\ : Odrv4
    port map (
            O => \N__25708\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3982\ : InMux
    port map (
            O => \N__25703\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__3981\ : InMux
    port map (
            O => \N__25700\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__3980\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25693\
        );

    \I__3979\ : InMux
    port map (
            O => \N__25696\,
            I => \N__25690\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__25693\,
            I => \N__25687\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__25690\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__25687\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3975\ : InMux
    port map (
            O => \N__25682\,
            I => \N__25678\
        );

    \I__3974\ : InMux
    port map (
            O => \N__25681\,
            I => \N__25674\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__25678\,
            I => \N__25671\
        );

    \I__3972\ : InMux
    port map (
            O => \N__25677\,
            I => \N__25668\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__25674\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3970\ : Odrv4
    port map (
            O => \N__25671\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__25668\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3968\ : InMux
    port map (
            O => \N__25661\,
            I => \bfn_11_6_0_\
        );

    \I__3967\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25654\
        );

    \I__3966\ : InMux
    port map (
            O => \N__25657\,
            I => \N__25651\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__25654\,
            I => \N__25648\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__25651\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3963\ : Odrv4
    port map (
            O => \N__25648\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3962\ : InMux
    port map (
            O => \N__25643\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__3961\ : InMux
    port map (
            O => \N__25640\,
            I => \N__25636\
        );

    \I__3960\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25633\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__25636\,
            I => \N__25630\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__25633\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__25630\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3956\ : InMux
    port map (
            O => \N__25625\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__3955\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25618\
        );

    \I__3954\ : InMux
    port map (
            O => \N__25621\,
            I => \N__25615\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__25618\,
            I => \N__25612\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__25615\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3951\ : Odrv12
    port map (
            O => \N__25612\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3950\ : InMux
    port map (
            O => \N__25607\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__3949\ : InMux
    port map (
            O => \N__25604\,
            I => \N__25600\
        );

    \I__3948\ : InMux
    port map (
            O => \N__25603\,
            I => \N__25597\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__25600\,
            I => \N__25594\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__25597\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3945\ : Odrv12
    port map (
            O => \N__25594\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3944\ : InMux
    port map (
            O => \N__25589\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__3943\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25582\
        );

    \I__3942\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25579\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__25582\,
            I => \N__25576\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__25579\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__25576\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3938\ : InMux
    port map (
            O => \N__25571\,
            I => \bfn_10_25_0_\
        );

    \I__3937\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25564\
        );

    \I__3936\ : InMux
    port map (
            O => \N__25567\,
            I => \N__25561\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__25564\,
            I => \N__25558\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__25561\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3933\ : Odrv4
    port map (
            O => \N__25558\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25553\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__3931\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25546\
        );

    \I__3930\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25543\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__25546\,
            I => \N__25540\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__25543\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__25540\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3926\ : InMux
    port map (
            O => \N__25535\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__3925\ : InMux
    port map (
            O => \N__25532\,
            I => \N__25528\
        );

    \I__3924\ : InMux
    port map (
            O => \N__25531\,
            I => \N__25525\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__25528\,
            I => \N__25522\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__25525\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__25522\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3920\ : InMux
    port map (
            O => \N__25517\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__3919\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25511\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__25511\,
            I => \phase_controller_inst2.stoper_hc.un6_running_19\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__25508\,
            I => \N__25505\
        );

    \I__3916\ : InMux
    port map (
            O => \N__25505\,
            I => \N__25502\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__25502\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\
        );

    \I__3914\ : InMux
    port map (
            O => \N__25499\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_19\
        );

    \I__3913\ : CascadeMux
    port map (
            O => \N__25496\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__3912\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25490\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__25490\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__3910\ : InMux
    port map (
            O => \N__25487\,
            I => \N__25483\
        );

    \I__3909\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25480\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__25483\,
            I => \N__25477\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__25480\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3906\ : Odrv4
    port map (
            O => \N__25477\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3905\ : InMux
    port map (
            O => \N__25472\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__25469\,
            I => \N__25466\
        );

    \I__3903\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__25463\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21\
        );

    \I__3901\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25456\
        );

    \I__3900\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25453\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__25456\,
            I => \N__25450\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__25453\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3897\ : Odrv4
    port map (
            O => \N__25450\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3896\ : InMux
    port map (
            O => \N__25445\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__3895\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25438\
        );

    \I__3894\ : InMux
    port map (
            O => \N__25441\,
            I => \N__25435\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__25438\,
            I => \N__25432\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__25435\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3891\ : Odrv4
    port map (
            O => \N__25432\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3890\ : InMux
    port map (
            O => \N__25427\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__3889\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25421\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__25421\,
            I => \phase_controller_inst2.stoper_hc.un6_running_11\
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__25418\,
            I => \N__25415\
        );

    \I__3886\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25412\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__25412\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__3884\ : CascadeMux
    port map (
            O => \N__25409\,
            I => \N__25406\
        );

    \I__3883\ : InMux
    port map (
            O => \N__25406\,
            I => \N__25403\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__25403\,
            I => \phase_controller_inst2.stoper_hc.un6_running_12\
        );

    \I__3881\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25397\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__25397\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__3879\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25391\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__25391\,
            I => \phase_controller_inst2.stoper_hc.un6_running_13\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__25388\,
            I => \N__25385\
        );

    \I__3876\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25382\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__25382\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__3874\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25376\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__25376\,
            I => \phase_controller_inst2.stoper_hc.un6_running_14\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__25373\,
            I => \N__25370\
        );

    \I__3871\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25367\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__25367\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__3869\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25361\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__25361\,
            I => \phase_controller_inst2.stoper_hc.un6_running_15\
        );

    \I__3867\ : CascadeMux
    port map (
            O => \N__25358\,
            I => \N__25355\
        );

    \I__3866\ : InMux
    port map (
            O => \N__25355\,
            I => \N__25352\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__25352\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__3864\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25346\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__25346\,
            I => \phase_controller_inst2.stoper_hc.un6_running_16\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__25343\,
            I => \N__25340\
        );

    \I__3861\ : InMux
    port map (
            O => \N__25340\,
            I => \N__25337\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__25337\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__25334\,
            I => \N__25331\
        );

    \I__3858\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25328\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__25328\,
            I => \phase_controller_inst2.stoper_hc.un6_running_17\
        );

    \I__3856\ : InMux
    port map (
            O => \N__25325\,
            I => \N__25322\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__25322\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\
        );

    \I__3854\ : InMux
    port map (
            O => \N__25319\,
            I => \N__25316\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__25316\,
            I => \phase_controller_inst2.stoper_hc.un6_running_18\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__25313\,
            I => \N__25310\
        );

    \I__3851\ : InMux
    port map (
            O => \N__25310\,
            I => \N__25307\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__25307\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\
        );

    \I__3849\ : InMux
    port map (
            O => \N__25304\,
            I => \N__25301\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__25301\,
            I => \N__25298\
        );

    \I__3847\ : Odrv4
    port map (
            O => \N__25298\,
            I => \phase_controller_inst2.stoper_hc.un6_running_3\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__25295\,
            I => \N__25292\
        );

    \I__3845\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25289\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__25289\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25286\,
            I => \N__25283\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__25283\,
            I => \N__25280\
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__25280\,
            I => \phase_controller_inst2.stoper_hc.un6_running_4\
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__25277\,
            I => \N__25274\
        );

    \I__3839\ : InMux
    port map (
            O => \N__25274\,
            I => \N__25271\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__25271\,
            I => \N__25268\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__25268\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__3836\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25262\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__25262\,
            I => \N__25259\
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__25259\,
            I => \phase_controller_inst2.stoper_hc.un6_running_5\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__25256\,
            I => \N__25253\
        );

    \I__3832\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25250\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__25250\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__3830\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25244\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__25244\,
            I => \N__25241\
        );

    \I__3828\ : Odrv4
    port map (
            O => \N__25241\,
            I => \phase_controller_inst2.stoper_hc.un6_running_6\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__25238\,
            I => \N__25235\
        );

    \I__3826\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25232\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__25232\,
            I => \N__25229\
        );

    \I__3824\ : Odrv4
    port map (
            O => \N__25229\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__3823\ : InMux
    port map (
            O => \N__25226\,
            I => \N__25223\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__25223\,
            I => \N__25220\
        );

    \I__3821\ : Odrv4
    port map (
            O => \N__25220\,
            I => \phase_controller_inst2.stoper_hc.un6_running_7\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__25217\,
            I => \N__25214\
        );

    \I__3819\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25211\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__25211\,
            I => \N__25208\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__25208\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__25205\,
            I => \N__25202\
        );

    \I__3815\ : InMux
    port map (
            O => \N__25202\,
            I => \N__25199\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__25199\,
            I => \N__25196\
        );

    \I__3813\ : Odrv4
    port map (
            O => \N__25196\,
            I => \phase_controller_inst2.stoper_hc.un6_running_8\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25190\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__25190\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25187\,
            I => \N__25184\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__25184\,
            I => \N__25181\
        );

    \I__3808\ : Span4Mux_v
    port map (
            O => \N__25181\,
            I => \N__25178\
        );

    \I__3807\ : Span4Mux_h
    port map (
            O => \N__25178\,
            I => \N__25175\
        );

    \I__3806\ : Odrv4
    port map (
            O => \N__25175\,
            I => \phase_controller_inst2.stoper_hc.un6_running_9\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__25172\,
            I => \N__25169\
        );

    \I__3804\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25166\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__25166\,
            I => \N__25163\
        );

    \I__3802\ : Odrv4
    port map (
            O => \N__25163\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__3801\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25157\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__25157\,
            I => \phase_controller_inst2.stoper_hc.un6_running_10\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__25154\,
            I => \N__25151\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25148\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__25148\,
            I => \N__25145\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__25145\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__3795\ : InMux
    port map (
            O => \N__25142\,
            I => \N__25139\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__25139\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15\
        );

    \I__3793\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25132\
        );

    \I__3792\ : InMux
    port map (
            O => \N__25135\,
            I => \N__25129\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__25132\,
            I => \elapsed_time_ns_1_RNI0AND11_0_28\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__25129\,
            I => \elapsed_time_ns_1_RNI0AND11_0_28\
        );

    \I__3789\ : InMux
    port map (
            O => \N__25124\,
            I => \N__25121\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__25121\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15\
        );

    \I__3787\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25112\
        );

    \I__3786\ : InMux
    port map (
            O => \N__25117\,
            I => \N__25112\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__25112\,
            I => \elapsed_time_ns_1_RNI1BND11_0_29\
        );

    \I__3784\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25105\
        );

    \I__3783\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25102\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__25105\,
            I => \elapsed_time_ns_1_RNIO1ND11_0_20\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__25102\,
            I => \elapsed_time_ns_1_RNIO1ND11_0_20\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__25097\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_\
        );

    \I__3779\ : InMux
    port map (
            O => \N__25094\,
            I => \N__25088\
        );

    \I__3778\ : InMux
    port map (
            O => \N__25093\,
            I => \N__25088\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__25088\,
            I => \elapsed_time_ns_1_RNIV8ND11_0_27\
        );

    \I__3776\ : CascadeMux
    port map (
            O => \N__25085\,
            I => \N__25082\
        );

    \I__3775\ : InMux
    port map (
            O => \N__25082\,
            I => \N__25079\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__3773\ : Odrv4
    port map (
            O => \N__25076\,
            I => \phase_controller_inst2.stoper_hc.un6_running_1\
        );

    \I__3772\ : InMux
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__25070\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__3770\ : InMux
    port map (
            O => \N__25067\,
            I => \N__25064\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__25064\,
            I => \N__25061\
        );

    \I__3768\ : Odrv4
    port map (
            O => \N__25061\,
            I => \phase_controller_inst2.stoper_hc.un6_running_2\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__25058\,
            I => \N__25055\
        );

    \I__3766\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__25049\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__25046\,
            I => \N__25043\
        );

    \I__3762\ : InMux
    port map (
            O => \N__25043\,
            I => \N__25039\
        );

    \I__3761\ : InMux
    port map (
            O => \N__25042\,
            I => \N__25035\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__25039\,
            I => \N__25032\
        );

    \I__3759\ : InMux
    port map (
            O => \N__25038\,
            I => \N__25028\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__25035\,
            I => \N__25023\
        );

    \I__3757\ : Span4Mux_v
    port map (
            O => \N__25032\,
            I => \N__25023\
        );

    \I__3756\ : InMux
    port map (
            O => \N__25031\,
            I => \N__25020\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__25028\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10\
        );

    \I__3754\ : Odrv4
    port map (
            O => \N__25023\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__25020\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10\
        );

    \I__3752\ : InMux
    port map (
            O => \N__25013\,
            I => \N__25010\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__25010\,
            I => \elapsed_time_ns_1_RNIP2ND11_0_21\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__25007\,
            I => \elapsed_time_ns_1_RNIP2ND11_0_21_cascade_\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__25004\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_\
        );

    \I__3748\ : InMux
    port map (
            O => \N__25001\,
            I => \N__24995\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24995\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__24995\,
            I => \elapsed_time_ns_1_RNIU7ND11_0_26\
        );

    \I__3745\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__24989\,
            I => \elapsed_time_ns_1_RNIR4ND11_0_23\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__24986\,
            I => \elapsed_time_ns_1_RNIR4ND11_0_23_cascade_\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__24983\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__24980\,
            I => \elapsed_time_ns_1_RNIP1MD11_0_12_cascade_\
        );

    \I__3740\ : InMux
    port map (
            O => \N__24977\,
            I => \N__24972\
        );

    \I__3739\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24969\
        );

    \I__3738\ : InMux
    port map (
            O => \N__24975\,
            I => \N__24966\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__24972\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__24969\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__24966\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\
        );

    \I__3734\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24954\
        );

    \I__3733\ : InMux
    port map (
            O => \N__24958\,
            I => \N__24949\
        );

    \I__3732\ : InMux
    port map (
            O => \N__24957\,
            I => \N__24949\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__24954\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__24949\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__24944\,
            I => \N__24940\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__24943\,
            I => \N__24936\
        );

    \I__3727\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24933\
        );

    \I__3726\ : InMux
    port map (
            O => \N__24939\,
            I => \N__24928\
        );

    \I__3725\ : InMux
    port map (
            O => \N__24936\,
            I => \N__24928\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__24933\,
            I => \N__24925\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__24928\,
            I => \N__24922\
        );

    \I__3722\ : Span4Mux_h
    port map (
            O => \N__24925\,
            I => \N__24919\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__24922\,
            I => \phase_controller_inst1.stoper_hc.N_337\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__24919\,
            I => \phase_controller_inst1.stoper_hc.N_337\
        );

    \I__3719\ : InMux
    port map (
            O => \N__24914\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__24911\,
            I => \N__24908\
        );

    \I__3717\ : InMux
    port map (
            O => \N__24908\,
            I => \N__24905\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__24905\,
            I => \N__24902\
        );

    \I__3715\ : Odrv4
    port map (
            O => \N__24902\,
            I => \current_shift_inst.PI_CTRL.integrator_i_29\
        );

    \I__3714\ : InMux
    port map (
            O => \N__24899\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\
        );

    \I__3713\ : InMux
    port map (
            O => \N__24896\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\
        );

    \I__3712\ : InMux
    port map (
            O => \N__24893\,
            I => \bfn_10_17_0_\
        );

    \I__3711\ : InMux
    port map (
            O => \N__24890\,
            I => \N__24887\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__24887\,
            I => \current_shift_inst.PI_CTRL.integrator_i_23\
        );

    \I__3709\ : InMux
    port map (
            O => \N__24884\,
            I => \N__24875\
        );

    \I__3708\ : InMux
    port map (
            O => \N__24883\,
            I => \N__24875\
        );

    \I__3707\ : InMux
    port map (
            O => \N__24882\,
            I => \N__24872\
        );

    \I__3706\ : InMux
    port map (
            O => \N__24881\,
            I => \N__24869\
        );

    \I__3705\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24866\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__24875\,
            I => \N__24863\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__24872\,
            I => \N__24860\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__24869\,
            I => \N__24855\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__24866\,
            I => \N__24855\
        );

    \I__3700\ : Span4Mux_h
    port map (
            O => \N__24863\,
            I => \N__24852\
        );

    \I__3699\ : Span4Mux_h
    port map (
            O => \N__24860\,
            I => \N__24847\
        );

    \I__3698\ : Span4Mux_h
    port map (
            O => \N__24855\,
            I => \N__24847\
        );

    \I__3697\ : Odrv4
    port map (
            O => \N__24852\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__24847\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3695\ : CascadeMux
    port map (
            O => \N__24842\,
            I => \N__24839\
        );

    \I__3694\ : InMux
    port map (
            O => \N__24839\,
            I => \N__24836\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__24836\,
            I => \N__24833\
        );

    \I__3692\ : Span4Mux_h
    port map (
            O => \N__24833\,
            I => \N__24830\
        );

    \I__3691\ : Odrv4
    port map (
            O => \N__24830\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\
        );

    \I__3690\ : InMux
    port map (
            O => \N__24827\,
            I => \N__24823\
        );

    \I__3689\ : InMux
    port map (
            O => \N__24826\,
            I => \N__24819\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__24823\,
            I => \N__24816\
        );

    \I__3687\ : InMux
    port map (
            O => \N__24822\,
            I => \N__24813\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__24819\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__3685\ : Odrv12
    port map (
            O => \N__24816\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__24813\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__24806\,
            I => \N__24803\
        );

    \I__3682\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24800\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__24800\,
            I => \N__24797\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__24797\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__24794\,
            I => \N__24791\
        );

    \I__3678\ : InMux
    port map (
            O => \N__24791\,
            I => \N__24788\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__24788\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\
        );

    \I__3676\ : InMux
    port map (
            O => \N__24785\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\
        );

    \I__3675\ : InMux
    port map (
            O => \N__24782\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\
        );

    \I__3674\ : InMux
    port map (
            O => \N__24779\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\
        );

    \I__3673\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24773\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__24773\,
            I => \N__24770\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__24770\,
            I => \N__24767\
        );

    \I__3670\ : Odrv4
    port map (
            O => \N__24767\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__3669\ : InMux
    port map (
            O => \N__24764\,
            I => \bfn_10_16_0_\
        );

    \I__3668\ : InMux
    port map (
            O => \N__24761\,
            I => \N__24758\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__24758\,
            I => \N__24755\
        );

    \I__3666\ : Span4Mux_h
    port map (
            O => \N__24755\,
            I => \N__24752\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__24752\,
            I => \current_shift_inst.PI_CTRL.integrator_i_24\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__24749\,
            I => \N__24746\
        );

    \I__3663\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24743\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__24743\,
            I => \N__24740\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__24740\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\
        );

    \I__3660\ : CascadeMux
    port map (
            O => \N__24737\,
            I => \N__24734\
        );

    \I__3659\ : InMux
    port map (
            O => \N__24734\,
            I => \N__24731\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__24731\,
            I => \N__24728\
        );

    \I__3657\ : Span4Mux_v
    port map (
            O => \N__24728\,
            I => \N__24725\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__24725\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__3655\ : InMux
    port map (
            O => \N__24722\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\
        );

    \I__3654\ : InMux
    port map (
            O => \N__24719\,
            I => \N__24716\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__24716\,
            I => \N__24713\
        );

    \I__3652\ : Span4Mux_v
    port map (
            O => \N__24713\,
            I => \N__24710\
        );

    \I__3651\ : Odrv4
    port map (
            O => \N__24710\,
            I => \current_shift_inst.PI_CTRL.integrator_i_25\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__24707\,
            I => \N__24704\
        );

    \I__3649\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24701\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__24701\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\
        );

    \I__3647\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24695\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__24695\,
            I => \N__24692\
        );

    \I__3645\ : Span4Mux_v
    port map (
            O => \N__24692\,
            I => \N__24689\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__24689\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__3643\ : InMux
    port map (
            O => \N__24686\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\
        );

    \I__3642\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24680\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__24680\,
            I => \N__24677\
        );

    \I__3640\ : Span12Mux_h
    port map (
            O => \N__24677\,
            I => \N__24674\
        );

    \I__3639\ : Odrv12
    port map (
            O => \N__24674\,
            I => \current_shift_inst.PI_CTRL.integrator_i_26\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__24671\,
            I => \N__24668\
        );

    \I__3637\ : InMux
    port map (
            O => \N__24668\,
            I => \N__24665\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__24665\,
            I => \N__24662\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__24662\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__24659\,
            I => \N__24656\
        );

    \I__3633\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24653\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__24653\,
            I => \N__24650\
        );

    \I__3631\ : Span4Mux_v
    port map (
            O => \N__24650\,
            I => \N__24647\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__24647\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__3629\ : InMux
    port map (
            O => \N__24644\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\
        );

    \I__3628\ : CascadeMux
    port map (
            O => \N__24641\,
            I => \N__24638\
        );

    \I__3627\ : InMux
    port map (
            O => \N__24638\,
            I => \N__24635\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__24635\,
            I => \N__24632\
        );

    \I__3625\ : Span4Mux_h
    port map (
            O => \N__24632\,
            I => \N__24629\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__24629\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__24626\,
            I => \N__24623\
        );

    \I__3622\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24620\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__3620\ : Odrv12
    port map (
            O => \N__24617\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__3619\ : InMux
    port map (
            O => \N__24614\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\
        );

    \I__3618\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__24608\,
            I => \N__24605\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__24605\,
            I => \current_shift_inst.PI_CTRL.integrator_i_12\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__24602\,
            I => \N__24599\
        );

    \I__3614\ : InMux
    port map (
            O => \N__24599\,
            I => \N__24596\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__24596\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\
        );

    \I__3612\ : InMux
    port map (
            O => \N__24593\,
            I => \N__24590\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__24590\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__3610\ : InMux
    port map (
            O => \N__24587\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\
        );

    \I__3609\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__24581\,
            I => \N__24578\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__24578\,
            I => \current_shift_inst.PI_CTRL.integrator_i_13\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__24575\,
            I => \N__24572\
        );

    \I__3605\ : InMux
    port map (
            O => \N__24572\,
            I => \N__24569\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__24569\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\
        );

    \I__3603\ : InMux
    port map (
            O => \N__24566\,
            I => \N__24563\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__24563\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__3601\ : InMux
    port map (
            O => \N__24560\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__24557\,
            I => \N__24554\
        );

    \I__3599\ : InMux
    port map (
            O => \N__24554\,
            I => \N__24551\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__24551\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\
        );

    \I__3597\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24545\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__24545\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__3595\ : InMux
    port map (
            O => \N__24542\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\
        );

    \I__3594\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__24536\,
            I => \N__24533\
        );

    \I__3592\ : Span4Mux_h
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__24530\,
            I => \current_shift_inst.PI_CTRL.integrator_i_15\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__24527\,
            I => \N__24524\
        );

    \I__3589\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24521\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__24521\,
            I => \N__24518\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__24518\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__24515\,
            I => \N__24512\
        );

    \I__3585\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24509\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__24509\,
            I => \N__24506\
        );

    \I__3583\ : Span4Mux_v
    port map (
            O => \N__24506\,
            I => \N__24503\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__24503\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__3581\ : InMux
    port map (
            O => \N__24500\,
            I => \bfn_10_15_0_\
        );

    \I__3580\ : InMux
    port map (
            O => \N__24497\,
            I => \N__24494\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__24494\,
            I => \N__24491\
        );

    \I__3578\ : Span4Mux_h
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__24488\,
            I => \current_shift_inst.PI_CTRL.integrator_i_16\
        );

    \I__3576\ : CascadeMux
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__3575\ : InMux
    port map (
            O => \N__24482\,
            I => \N__24479\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__24479\,
            I => \N__24476\
        );

    \I__3573\ : Span4Mux_h
    port map (
            O => \N__24476\,
            I => \N__24473\
        );

    \I__3572\ : Odrv4
    port map (
            O => \N__24473\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\
        );

    \I__3571\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24467\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__24467\,
            I => \N__24464\
        );

    \I__3569\ : Span4Mux_v
    port map (
            O => \N__24464\,
            I => \N__24461\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__24461\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__3567\ : InMux
    port map (
            O => \N__24458\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\
        );

    \I__3566\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24452\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__24452\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__3563\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24443\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__24443\,
            I => \current_shift_inst.PI_CTRL.integrator_i_17\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__24440\,
            I => \N__24437\
        );

    \I__3560\ : InMux
    port map (
            O => \N__24437\,
            I => \N__24434\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__24434\,
            I => \N__24431\
        );

    \I__3558\ : Span4Mux_h
    port map (
            O => \N__24431\,
            I => \N__24428\
        );

    \I__3557\ : Span4Mux_h
    port map (
            O => \N__24428\,
            I => \N__24425\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__24425\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__3555\ : InMux
    port map (
            O => \N__24422\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\
        );

    \I__3554\ : InMux
    port map (
            O => \N__24419\,
            I => \N__24416\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__24416\,
            I => \N__24413\
        );

    \I__3552\ : Span4Mux_v
    port map (
            O => \N__24413\,
            I => \N__24410\
        );

    \I__3551\ : Odrv4
    port map (
            O => \N__24410\,
            I => \current_shift_inst.PI_CTRL.integrator_i_18\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__24407\,
            I => \N__24404\
        );

    \I__3549\ : InMux
    port map (
            O => \N__24404\,
            I => \N__24401\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__24401\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\
        );

    \I__3547\ : InMux
    port map (
            O => \N__24398\,
            I => \N__24395\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__3545\ : Span4Mux_h
    port map (
            O => \N__24392\,
            I => \N__24389\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__24389\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__3543\ : InMux
    port map (
            O => \N__24386\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__24383\,
            I => \N__24380\
        );

    \I__3541\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24377\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__24377\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\
        );

    \I__3539\ : InMux
    port map (
            O => \N__24374\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\
        );

    \I__3538\ : InMux
    port map (
            O => \N__24371\,
            I => \N__24368\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__24368\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__3536\ : InMux
    port map (
            O => \N__24365\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24359\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24356\
        );

    \I__3533\ : Span4Mux_v
    port map (
            O => \N__24356\,
            I => \N__24353\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__24353\,
            I => \current_shift_inst.PI_CTRL.integrator_i_5\
        );

    \I__3531\ : InMux
    port map (
            O => \N__24350\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\
        );

    \I__3530\ : InMux
    port map (
            O => \N__24347\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\
        );

    \I__3529\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24341\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__24341\,
            I => \N__24338\
        );

    \I__3527\ : Odrv4
    port map (
            O => \N__24338\,
            I => \current_shift_inst.PI_CTRL.integrator_i_7\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__24335\,
            I => \N__24332\
        );

    \I__3525\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24326\
        );

    \I__3523\ : Span4Mux_h
    port map (
            O => \N__24326\,
            I => \N__24323\
        );

    \I__3522\ : Odrv4
    port map (
            O => \N__24323\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\
        );

    \I__3521\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24317\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__24317\,
            I => \N__24314\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__24314\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__3518\ : InMux
    port map (
            O => \N__24311\,
            I => \bfn_10_14_0_\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24305\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24302\
        );

    \I__3515\ : Odrv4
    port map (
            O => \N__24302\,
            I => \current_shift_inst.PI_CTRL.integrator_i_8\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__24299\,
            I => \N__24296\
        );

    \I__3513\ : InMux
    port map (
            O => \N__24296\,
            I => \N__24293\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__24293\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\
        );

    \I__3511\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__24287\,
            I => \N__24284\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__24284\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__3508\ : InMux
    port map (
            O => \N__24281\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\
        );

    \I__3507\ : InMux
    port map (
            O => \N__24278\,
            I => \N__24275\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__24275\,
            I => \N__24272\
        );

    \I__3505\ : Span4Mux_v
    port map (
            O => \N__24272\,
            I => \N__24269\
        );

    \I__3504\ : Odrv4
    port map (
            O => \N__24269\,
            I => \current_shift_inst.PI_CTRL.integrator_i_9\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__24266\,
            I => \N__24263\
        );

    \I__3502\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24260\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__24260\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__24257\,
            I => \N__24254\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24251\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__3497\ : Odrv4
    port map (
            O => \N__24248\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24245\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__24242\,
            I => \N__24239\
        );

    \I__3494\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24236\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__24236\,
            I => \N__24233\
        );

    \I__3492\ : Odrv4
    port map (
            O => \N__24233\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24230\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24227\,
            I => \N__24224\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__24224\,
            I => \N__24221\
        );

    \I__3488\ : Odrv12
    port map (
            O => \N__24221\,
            I => \current_shift_inst.PI_CTRL.integrator_i_11\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__24218\,
            I => \N__24215\
        );

    \I__3486\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24212\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__24212\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__24203\,
            I => \N__24200\
        );

    \I__3481\ : Odrv4
    port map (
            O => \N__24200\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__3480\ : InMux
    port map (
            O => \N__24197\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__3478\ : InMux
    port map (
            O => \N__24191\,
            I => \N__24187\
        );

    \I__3477\ : InMux
    port map (
            O => \N__24190\,
            I => \N__24184\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__24187\,
            I => \N__24181\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__24184\,
            I => \N__24176\
        );

    \I__3474\ : Span4Mux_h
    port map (
            O => \N__24181\,
            I => \N__24173\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24180\,
            I => \N__24168\
        );

    \I__3472\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24168\
        );

    \I__3471\ : Span4Mux_h
    port map (
            O => \N__24176\,
            I => \N__24162\
        );

    \I__3470\ : Span4Mux_h
    port map (
            O => \N__24173\,
            I => \N__24162\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__24168\,
            I => \N__24159\
        );

    \I__3468\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24156\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__24162\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__24159\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__24156\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3464\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24145\
        );

    \I__3463\ : InMux
    port map (
            O => \N__24148\,
            I => \N__24142\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__24145\,
            I => \N__24139\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__24142\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__24139\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__24134\,
            I => \N__24131\
        );

    \I__3458\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24128\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__24128\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\
        );

    \I__3456\ : CascadeMux
    port map (
            O => \N__24125\,
            I => \N__24121\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__24124\,
            I => \N__24118\
        );

    \I__3454\ : InMux
    port map (
            O => \N__24121\,
            I => \N__24115\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24112\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__24115\,
            I => \N__24108\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__24112\,
            I => \N__24105\
        );

    \I__3450\ : InMux
    port map (
            O => \N__24111\,
            I => \N__24102\
        );

    \I__3449\ : Span12Mux_s10_h
    port map (
            O => \N__24108\,
            I => \N__24099\
        );

    \I__3448\ : Span4Mux_v
    port map (
            O => \N__24105\,
            I => \N__24094\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__24102\,
            I => \N__24094\
        );

    \I__3446\ : Odrv12
    port map (
            O => \N__24099\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__24094\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3444\ : InMux
    port map (
            O => \N__24089\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\
        );

    \I__3443\ : InMux
    port map (
            O => \N__24086\,
            I => \N__24083\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__24083\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\
        );

    \I__3441\ : InMux
    port map (
            O => \N__24080\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\
        );

    \I__3440\ : InMux
    port map (
            O => \N__24077\,
            I => \N__24074\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__24074\,
            I => \N__24071\
        );

    \I__3438\ : Span4Mux_h
    port map (
            O => \N__24071\,
            I => \N__24068\
        );

    \I__3437\ : Span4Mux_h
    port map (
            O => \N__24068\,
            I => \N__24065\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__24065\,
            I => \current_shift_inst.PI_CTRL.integrator_i_2\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__24062\,
            I => \N__24059\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24059\,
            I => \N__24056\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__24056\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__24053\,
            I => \N__24050\
        );

    \I__3431\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24045\
        );

    \I__3430\ : InMux
    port map (
            O => \N__24049\,
            I => \N__24042\
        );

    \I__3429\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24039\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__24045\,
            I => \N__24035\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__24042\,
            I => \N__24032\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__24039\,
            I => \N__24029\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24026\
        );

    \I__3424\ : Span4Mux_h
    port map (
            O => \N__24035\,
            I => \N__24023\
        );

    \I__3423\ : Span4Mux_h
    port map (
            O => \N__24032\,
            I => \N__24020\
        );

    \I__3422\ : Span4Mux_v
    port map (
            O => \N__24029\,
            I => \N__24017\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__24026\,
            I => \N__24010\
        );

    \I__3420\ : Span4Mux_h
    port map (
            O => \N__24023\,
            I => \N__24010\
        );

    \I__3419\ : Span4Mux_h
    port map (
            O => \N__24020\,
            I => \N__24010\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__24017\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__24010\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__3416\ : InMux
    port map (
            O => \N__24005\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\
        );

    \I__3415\ : InMux
    port map (
            O => \N__24002\,
            I => \N__23999\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__23999\,
            I => \N__23996\
        );

    \I__3413\ : Odrv12
    port map (
            O => \N__23996\,
            I => \current_shift_inst.PI_CTRL.integrator_i_3\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__23993\,
            I => \N__23990\
        );

    \I__3411\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23987\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__23987\,
            I => \N__23984\
        );

    \I__3409\ : Odrv4
    port map (
            O => \N__23984\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__23981\,
            I => \N__23977\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__23980\,
            I => \N__23974\
        );

    \I__3406\ : InMux
    port map (
            O => \N__23977\,
            I => \N__23970\
        );

    \I__3405\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23966\
        );

    \I__3404\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23963\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__23970\,
            I => \N__23960\
        );

    \I__3402\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23956\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__23966\,
            I => \N__23951\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__23963\,
            I => \N__23951\
        );

    \I__3399\ : Span4Mux_v
    port map (
            O => \N__23960\,
            I => \N__23948\
        );

    \I__3398\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23945\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__23956\,
            I => \N__23938\
        );

    \I__3396\ : Span4Mux_h
    port map (
            O => \N__23951\,
            I => \N__23938\
        );

    \I__3395\ : Span4Mux_h
    port map (
            O => \N__23948\,
            I => \N__23938\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__23945\,
            I => \N__23935\
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__23938\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3392\ : Odrv4
    port map (
            O => \N__23935\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3391\ : InMux
    port map (
            O => \N__23930\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\
        );

    \I__3390\ : InMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__23924\,
            I => \current_shift_inst.PI_CTRL.integrator_i_4\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__23921\,
            I => \N__23918\
        );

    \I__3387\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23915\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__23915\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__23912\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__3384\ : InMux
    port map (
            O => \N__23909\,
            I => \N__23906\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__23906\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__23903\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__3381\ : InMux
    port map (
            O => \N__23900\,
            I => \N__23897\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__23897\,
            I => \N__23894\
        );

    \I__3379\ : Span4Mux_h
    port map (
            O => \N__23894\,
            I => \N__23891\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__23891\,
            I => \il_max_comp2_D1\
        );

    \I__3377\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__23885\,
            I => \il_min_comp1_D1\
        );

    \I__3375\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23875\
        );

    \I__3373\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23872\
        );

    \I__3372\ : Span4Mux_h
    port map (
            O => \N__23875\,
            I => \N__23869\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__23872\,
            I => \N__23861\
        );

    \I__3370\ : Span4Mux_h
    port map (
            O => \N__23869\,
            I => \N__23861\
        );

    \I__3369\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23856\
        );

    \I__3368\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23856\
        );

    \I__3367\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23853\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__23861\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__23856\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__23853\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3363\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23842\
        );

    \I__3362\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23839\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__23842\,
            I => \phase_controller_inst1.stoper_hc.N_287\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__23839\,
            I => \phase_controller_inst1.stoper_hc.N_287\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__23834\,
            I => \N__23830\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__23833\,
            I => \N__23824\
        );

    \I__3357\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23821\
        );

    \I__3356\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23818\
        );

    \I__3355\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23815\
        );

    \I__3354\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23810\
        );

    \I__3353\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23807\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__23821\,
            I => \N__23804\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__23818\,
            I => \N__23801\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__23815\,
            I => \N__23798\
        );

    \I__3349\ : InMux
    port map (
            O => \N__23814\,
            I => \N__23795\
        );

    \I__3348\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23792\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__23810\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__23807\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__23804\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__23801\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__3343\ : Odrv4
    port map (
            O => \N__23798\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__23795\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__23792\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23777\,
            I => \N__23773\
        );

    \I__3339\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23770\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__23773\,
            I => \N__23764\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__23770\,
            I => \N__23764\
        );

    \I__3336\ : InMux
    port map (
            O => \N__23769\,
            I => \N__23759\
        );

    \I__3335\ : Span4Mux_v
    port map (
            O => \N__23764\,
            I => \N__23756\
        );

    \I__3334\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23751\
        );

    \I__3333\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23751\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__23759\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18\
        );

    \I__3331\ : Odrv4
    port map (
            O => \N__23756\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__23751\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18\
        );

    \I__3329\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23739\
        );

    \I__3328\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23736\
        );

    \I__3327\ : InMux
    port map (
            O => \N__23742\,
            I => \N__23733\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__23739\,
            I => \N__23727\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__23736\,
            I => \N__23727\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__23733\,
            I => \N__23724\
        );

    \I__3323\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23721\
        );

    \I__3322\ : Odrv4
    port map (
            O => \N__23727\,
            I => \elapsed_time_ns_1_RNI40CED1_0_17\
        );

    \I__3321\ : Odrv4
    port map (
            O => \N__23724\,
            I => \elapsed_time_ns_1_RNI40CED1_0_17\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__23721\,
            I => \elapsed_time_ns_1_RNI40CED1_0_17\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__23714\,
            I => \N__23709\
        );

    \I__3318\ : InMux
    port map (
            O => \N__23713\,
            I => \N__23704\
        );

    \I__3317\ : InMux
    port map (
            O => \N__23712\,
            I => \N__23701\
        );

    \I__3316\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23696\
        );

    \I__3315\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23696\
        );

    \I__3314\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23693\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__23704\,
            I => \N__23690\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__23701\,
            I => \N__23685\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__23696\,
            I => \N__23685\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__23693\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__23690\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19\
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__23685\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19\
        );

    \I__3307\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23674\
        );

    \I__3306\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23671\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__23674\,
            I => \N__23666\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__23671\,
            I => \N__23666\
        );

    \I__3303\ : Span4Mux_v
    port map (
            O => \N__23666\,
            I => \N__23661\
        );

    \I__3302\ : InMux
    port map (
            O => \N__23665\,
            I => \N__23658\
        );

    \I__3301\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23655\
        );

    \I__3300\ : Span4Mux_h
    port map (
            O => \N__23661\,
            I => \N__23652\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__23658\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__23655\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__3297\ : Odrv4
    port map (
            O => \N__23652\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__3296\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23641\
        );

    \I__3295\ : InMux
    port map (
            O => \N__23644\,
            I => \N__23637\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__23641\,
            I => \N__23634\
        );

    \I__3293\ : InMux
    port map (
            O => \N__23640\,
            I => \N__23631\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__23637\,
            I => \N__23624\
        );

    \I__3291\ : Span4Mux_h
    port map (
            O => \N__23634\,
            I => \N__23624\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__23631\,
            I => \N__23624\
        );

    \I__3289\ : Span4Mux_h
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__3288\ : Span4Mux_v
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__23618\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__3286\ : IoInMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__23609\,
            I => s3_phy_c
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__23606\,
            I => \N__23602\
        );

    \I__3282\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23596\
        );

    \I__3281\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23593\
        );

    \I__3280\ : InMux
    port map (
            O => \N__23601\,
            I => \N__23590\
        );

    \I__3279\ : InMux
    port map (
            O => \N__23600\,
            I => \N__23585\
        );

    \I__3278\ : InMux
    port map (
            O => \N__23599\,
            I => \N__23585\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__23596\,
            I => \elapsed_time_ns_1_RNIL13KD1_0_9\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__23593\,
            I => \elapsed_time_ns_1_RNIL13KD1_0_9\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__23590\,
            I => \elapsed_time_ns_1_RNIL13KD1_0_9\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__23585\,
            I => \elapsed_time_ns_1_RNIL13KD1_0_9\
        );

    \I__3273\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__23573\,
            I => \N__23569\
        );

    \I__3271\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23566\
        );

    \I__3270\ : Span4Mux_v
    port map (
            O => \N__23569\,
            I => \N__23563\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__23566\,
            I => \N__23560\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__23563\,
            I => \phase_controller_inst1.stoper_hc.N_266_iZ0Z_1\
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__23560\,
            I => \phase_controller_inst1.stoper_hc.N_266_iZ0Z_1\
        );

    \I__3266\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23551\
        );

    \I__3265\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23546\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__23551\,
            I => \N__23543\
        );

    \I__3263\ : InMux
    port map (
            O => \N__23550\,
            I => \N__23538\
        );

    \I__3262\ : InMux
    port map (
            O => \N__23549\,
            I => \N__23538\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__23546\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16\
        );

    \I__3260\ : Odrv4
    port map (
            O => \N__23543\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__23538\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__23531\,
            I => \phase_controller_inst1.stoper_hc.N_325_cascade_\
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__23528\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__23525\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5_cascade_\
        );

    \I__3255\ : CascadeMux
    port map (
            O => \N__23522\,
            I => \N__23518\
        );

    \I__3254\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23515\
        );

    \I__3253\ : InMux
    port map (
            O => \N__23518\,
            I => \N__23512\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__23515\,
            I => \N__23508\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__23512\,
            I => \N__23505\
        );

    \I__3250\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23502\
        );

    \I__3249\ : Span4Mux_h
    port map (
            O => \N__23508\,
            I => \N__23495\
        );

    \I__3248\ : Span4Mux_h
    port map (
            O => \N__23505\,
            I => \N__23495\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__23502\,
            I => \N__23492\
        );

    \I__3246\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23487\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23487\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__23495\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__23492\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__23487\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3241\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23476\
        );

    \I__3240\ : InMux
    port map (
            O => \N__23479\,
            I => \N__23472\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__23476\,
            I => \N__23469\
        );

    \I__3238\ : InMux
    port map (
            O => \N__23475\,
            I => \N__23466\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__23472\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__23469\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__23466\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__3234\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23456\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__23456\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\
        );

    \I__3232\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23449\
        );

    \I__3231\ : InMux
    port map (
            O => \N__23452\,
            I => \N__23446\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__23449\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__23446\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__3228\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23438\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__23438\,
            I => \N__23435\
        );

    \I__3226\ : Odrv4
    port map (
            O => \N__23435\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__23432\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_\
        );

    \I__3224\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23424\
        );

    \I__3223\ : InMux
    port map (
            O => \N__23428\,
            I => \N__23421\
        );

    \I__3222\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23418\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__23424\,
            I => \N__23413\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__23421\,
            I => \N__23410\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__23418\,
            I => \N__23407\
        );

    \I__3218\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23402\
        );

    \I__3217\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23402\
        );

    \I__3216\ : Span4Mux_h
    port map (
            O => \N__23413\,
            I => \N__23397\
        );

    \I__3215\ : Span4Mux_h
    port map (
            O => \N__23410\,
            I => \N__23397\
        );

    \I__3214\ : Span4Mux_h
    port map (
            O => \N__23407\,
            I => \N__23392\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__23402\,
            I => \N__23392\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__23397\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__23392\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3210\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23383\
        );

    \I__3209\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23380\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__23383\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__23380\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__3206\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23371\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__23374\,
            I => \N__23368\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__23371\,
            I => \N__23365\
        );

    \I__3203\ : InMux
    port map (
            O => \N__23368\,
            I => \N__23362\
        );

    \I__3202\ : Span4Mux_v
    port map (
            O => \N__23365\,
            I => \N__23357\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__23362\,
            I => \N__23354\
        );

    \I__3200\ : InMux
    port map (
            O => \N__23361\,
            I => \N__23351\
        );

    \I__3199\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23348\
        );

    \I__3198\ : Span4Mux_h
    port map (
            O => \N__23357\,
            I => \N__23342\
        );

    \I__3197\ : Span4Mux_v
    port map (
            O => \N__23354\,
            I => \N__23342\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__23351\,
            I => \N__23339\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__23348\,
            I => \N__23336\
        );

    \I__3194\ : InMux
    port map (
            O => \N__23347\,
            I => \N__23333\
        );

    \I__3193\ : Odrv4
    port map (
            O => \N__23342\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__23339\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__23336\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__23333\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__23324\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_\
        );

    \I__3188\ : InMux
    port map (
            O => \N__23321\,
            I => \N__23318\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__23318\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\
        );

    \I__3186\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23311\
        );

    \I__3185\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23307\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__23311\,
            I => \N__23304\
        );

    \I__3183\ : InMux
    port map (
            O => \N__23310\,
            I => \N__23301\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__23307\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__3181\ : Odrv12
    port map (
            O => \N__23304\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__23301\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__23294\,
            I => \N__23291\
        );

    \I__3178\ : InMux
    port map (
            O => \N__23291\,
            I => \N__23286\
        );

    \I__3177\ : InMux
    port map (
            O => \N__23290\,
            I => \N__23283\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__23289\,
            I => \N__23280\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__23286\,
            I => \N__23276\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__23283\,
            I => \N__23273\
        );

    \I__3173\ : InMux
    port map (
            O => \N__23280\,
            I => \N__23270\
        );

    \I__3172\ : InMux
    port map (
            O => \N__23279\,
            I => \N__23267\
        );

    \I__3171\ : Span4Mux_h
    port map (
            O => \N__23276\,
            I => \N__23263\
        );

    \I__3170\ : Span4Mux_v
    port map (
            O => \N__23273\,
            I => \N__23256\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__23270\,
            I => \N__23256\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__23267\,
            I => \N__23256\
        );

    \I__3167\ : InMux
    port map (
            O => \N__23266\,
            I => \N__23253\
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__23263\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3165\ : Odrv4
    port map (
            O => \N__23256\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__23253\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__3162\ : InMux
    port map (
            O => \N__23243\,
            I => \N__23240\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__23240\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__23237\,
            I => \phase_controller_inst1.stoper_hc.N_275_cascade_\
        );

    \I__3159\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23230\
        );

    \I__3158\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23227\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__23230\,
            I => \N__23224\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__23227\,
            I => \N__23218\
        );

    \I__3155\ : Span4Mux_h
    port map (
            O => \N__23224\,
            I => \N__23215\
        );

    \I__3154\ : InMux
    port map (
            O => \N__23223\,
            I => \N__23212\
        );

    \I__3153\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23209\
        );

    \I__3152\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23206\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__23218\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__23215\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__23212\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__23209\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__23206\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3146\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23191\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23188\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__23191\,
            I => \N__23182\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__23188\,
            I => \N__23182\
        );

    \I__3142\ : InMux
    port map (
            O => \N__23187\,
            I => \N__23179\
        );

    \I__3141\ : Sp12to4
    port map (
            O => \N__23182\,
            I => \N__23176\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__23179\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__3139\ : Odrv12
    port map (
            O => \N__23176\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__3138\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23168\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23165\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__23165\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\
        );

    \I__3135\ : InMux
    port map (
            O => \N__23162\,
            I => \N__23159\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__23159\,
            I => \N__23156\
        );

    \I__3133\ : Span4Mux_v
    port map (
            O => \N__23156\,
            I => \N__23153\
        );

    \I__3132\ : Odrv4
    port map (
            O => \N__23153\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__3131\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23147\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__23147\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23140\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23135\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__23140\,
            I => \N__23132\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__23139\,
            I => \N__23129\
        );

    \I__3125\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23125\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__23135\,
            I => \N__23122\
        );

    \I__3123\ : Span4Mux_h
    port map (
            O => \N__23132\,
            I => \N__23119\
        );

    \I__3122\ : InMux
    port map (
            O => \N__23129\,
            I => \N__23116\
        );

    \I__3121\ : InMux
    port map (
            O => \N__23128\,
            I => \N__23113\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__23125\,
            I => \N__23110\
        );

    \I__3119\ : Odrv4
    port map (
            O => \N__23122\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__23119\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__23116\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__23113\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__23110\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__23099\,
            I => \N__23096\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23093\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__23093\,
            I => \N__23089\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23085\
        );

    \I__3110\ : Span4Mux_h
    port map (
            O => \N__23089\,
            I => \N__23082\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23079\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__23085\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__23082\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__23079\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__3105\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23069\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__23069\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__23066\,
            I => \N__23062\
        );

    \I__3102\ : InMux
    port map (
            O => \N__23065\,
            I => \N__23058\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23062\,
            I => \N__23055\
        );

    \I__3100\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23052\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__23058\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__23055\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__23052\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__3096\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23042\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__23042\,
            I => \N__23039\
        );

    \I__3094\ : Odrv4
    port map (
            O => \N__23039\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23033\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__23033\,
            I => \N__23028\
        );

    \I__3091\ : InMux
    port map (
            O => \N__23032\,
            I => \N__23025\
        );

    \I__3090\ : InMux
    port map (
            O => \N__23031\,
            I => \N__23022\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__23028\,
            I => \N__23017\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__23025\,
            I => \N__23017\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__23022\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__23017\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23012\,
            I => \N__23007\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23011\,
            I => \N__23004\
        );

    \I__3083\ : InMux
    port map (
            O => \N__23010\,
            I => \N__23001\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__23007\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__23004\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__23001\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__22994\,
            I => \N__22991\
        );

    \I__3078\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22986\
        );

    \I__3077\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22982\
        );

    \I__3076\ : InMux
    port map (
            O => \N__22989\,
            I => \N__22979\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__22986\,
            I => \N__22976\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__22985\,
            I => \N__22972\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__22982\,
            I => \N__22969\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__22979\,
            I => \N__22966\
        );

    \I__3071\ : Span4Mux_h
    port map (
            O => \N__22976\,
            I => \N__22963\
        );

    \I__3070\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22960\
        );

    \I__3069\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22957\
        );

    \I__3068\ : Span4Mux_v
    port map (
            O => \N__22969\,
            I => \N__22954\
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__22966\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__22963\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__22960\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__22957\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__22954\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3062\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22940\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__22940\,
            I => \N__22936\
        );

    \I__3060\ : InMux
    port map (
            O => \N__22939\,
            I => \N__22932\
        );

    \I__3059\ : Span4Mux_v
    port map (
            O => \N__22936\,
            I => \N__22929\
        );

    \I__3058\ : InMux
    port map (
            O => \N__22935\,
            I => \N__22926\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__22932\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__22929\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__22926\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__22919\,
            I => \N__22916\
        );

    \I__3053\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22913\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__22913\,
            I => \N__22910\
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__22910\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__22907\,
            I => \N__22903\
        );

    \I__3049\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22900\
        );

    \I__3048\ : InMux
    port map (
            O => \N__22903\,
            I => \N__22897\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__22900\,
            I => \N__22892\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__22897\,
            I => \N__22889\
        );

    \I__3045\ : InMux
    port map (
            O => \N__22896\,
            I => \N__22885\
        );

    \I__3044\ : InMux
    port map (
            O => \N__22895\,
            I => \N__22882\
        );

    \I__3043\ : Span4Mux_v
    port map (
            O => \N__22892\,
            I => \N__22879\
        );

    \I__3042\ : Span4Mux_v
    port map (
            O => \N__22889\,
            I => \N__22876\
        );

    \I__3041\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22873\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__22885\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__22882\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__22879\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3037\ : Odrv4
    port map (
            O => \N__22876\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__22873\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__22862\,
            I => \N__22858\
        );

    \I__3034\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22855\
        );

    \I__3033\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22852\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__22855\,
            I => \N__22849\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__22852\,
            I => \N__22846\
        );

    \I__3030\ : Span4Mux_v
    port map (
            O => \N__22849\,
            I => \N__22842\
        );

    \I__3029\ : Span4Mux_h
    port map (
            O => \N__22846\,
            I => \N__22839\
        );

    \I__3028\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22836\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__22842\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__22839\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__22836\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__3024\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22826\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__22823\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_8\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__22820\,
            I => \N__22817\
        );

    \I__3020\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22813\
        );

    \I__3019\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22809\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__22813\,
            I => \N__22806\
        );

    \I__3017\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22803\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__22809\,
            I => \N__22800\
        );

    \I__3015\ : Span4Mux_v
    port map (
            O => \N__22806\,
            I => \N__22797\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__22803\,
            I => \N__22794\
        );

    \I__3013\ : Odrv12
    port map (
            O => \N__22800\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__3012\ : Odrv4
    port map (
            O => \N__22797\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__22794\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__3010\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22784\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__22784\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\
        );

    \I__3008\ : InMux
    port map (
            O => \N__22781\,
            I => \N__22778\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__22778\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__3005\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22767\
        );

    \I__3004\ : InMux
    port map (
            O => \N__22771\,
            I => \N__22764\
        );

    \I__3003\ : InMux
    port map (
            O => \N__22770\,
            I => \N__22761\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__22767\,
            I => \N__22758\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__22764\,
            I => \N__22755\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__22761\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__2999\ : Odrv4
    port map (
            O => \N__22758\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__2998\ : Odrv12
    port map (
            O => \N__22755\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__2997\ : InMux
    port map (
            O => \N__22748\,
            I => \N__22745\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__22745\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\
        );

    \I__2995\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22738\
        );

    \I__2994\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22735\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__22738\,
            I => \N__22732\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22726\
        );

    \I__2991\ : Span4Mux_v
    port map (
            O => \N__22732\,
            I => \N__22723\
        );

    \I__2990\ : InMux
    port map (
            O => \N__22731\,
            I => \N__22720\
        );

    \I__2989\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22715\
        );

    \I__2988\ : InMux
    port map (
            O => \N__22729\,
            I => \N__22715\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__22726\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2986\ : Odrv4
    port map (
            O => \N__22723\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__22720\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__22715\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2983\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22702\
        );

    \I__2982\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22699\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__22702\,
            I => \N__22696\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__22699\,
            I => \N__22690\
        );

    \I__2979\ : Span4Mux_v
    port map (
            O => \N__22696\,
            I => \N__22690\
        );

    \I__2978\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22687\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__22690\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__22687\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__2975\ : InMux
    port map (
            O => \N__22682\,
            I => \N__22679\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__2973\ : Odrv4
    port map (
            O => \N__22676\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\
        );

    \I__2972\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22669\
        );

    \I__2971\ : InMux
    port map (
            O => \N__22672\,
            I => \N__22666\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__22669\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__22666\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__22661\,
            I => \N__22657\
        );

    \I__2967\ : InMux
    port map (
            O => \N__22660\,
            I => \N__22654\
        );

    \I__2966\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22651\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__22654\,
            I => \N__22645\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__22651\,
            I => \N__22642\
        );

    \I__2963\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22639\
        );

    \I__2962\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22633\
        );

    \I__2961\ : InMux
    port map (
            O => \N__22648\,
            I => \N__22633\
        );

    \I__2960\ : Span4Mux_h
    port map (
            O => \N__22645\,
            I => \N__22626\
        );

    \I__2959\ : Span4Mux_h
    port map (
            O => \N__22642\,
            I => \N__22626\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__22639\,
            I => \N__22626\
        );

    \I__2957\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22623\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__22633\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__22626\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__22623\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__22616\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_\
        );

    \I__2952\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22610\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__22610\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__22607\,
            I => \N__22604\
        );

    \I__2949\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22601\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22598\
        );

    \I__2947\ : Odrv12
    port map (
            O => \N__22598\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_7\
        );

    \I__2946\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22592\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__22592\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\
        );

    \I__2944\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22586\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__2942\ : Span4Mux_h
    port map (
            O => \N__22583\,
            I => \N__22580\
        );

    \I__2941\ : Odrv4
    port map (
            O => \N__22580\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\
        );

    \I__2940\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22574\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__22574\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_4\
        );

    \I__2938\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22568\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__22568\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_5\
        );

    \I__2936\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__22562\,
            I => \N__22559\
        );

    \I__2934\ : Span4Mux_v
    port map (
            O => \N__22559\,
            I => \N__22555\
        );

    \I__2933\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22551\
        );

    \I__2932\ : Span4Mux_h
    port map (
            O => \N__22555\,
            I => \N__22548\
        );

    \I__2931\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22545\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__22551\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__2929\ : Odrv4
    port map (
            O => \N__22548\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__22545\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__2927\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__22535\,
            I => \N__22532\
        );

    \I__2925\ : Odrv4
    port map (
            O => \N__22532\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\
        );

    \I__2924\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22526\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__22526\,
            I => \N__22522\
        );

    \I__2922\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22518\
        );

    \I__2921\ : Span4Mux_h
    port map (
            O => \N__22522\,
            I => \N__22515\
        );

    \I__2920\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22512\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__22518\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__2918\ : Odrv4
    port map (
            O => \N__22515\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__22512\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__22505\,
            I => \N__22502\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22493\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__22498\,
            I => \N__22490\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__22497\,
            I => \N__22487\
        );

    \I__2911\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22483\
        );

    \I__2910\ : Span4Mux_v
    port map (
            O => \N__22493\,
            I => \N__22480\
        );

    \I__2909\ : InMux
    port map (
            O => \N__22490\,
            I => \N__22475\
        );

    \I__2908\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22475\
        );

    \I__2907\ : InMux
    port map (
            O => \N__22486\,
            I => \N__22472\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__22483\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__22480\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__22475\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__22472\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2902\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22460\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__22460\,
            I => \N__22457\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__22457\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\
        );

    \I__2899\ : InMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__22451\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_6\
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__2896\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22441\
        );

    \I__2895\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22437\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__22441\,
            I => \N__22434\
        );

    \I__2893\ : InMux
    port map (
            O => \N__22440\,
            I => \N__22431\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__22437\,
            I => \N__22428\
        );

    \I__2891\ : Span4Mux_h
    port map (
            O => \N__22434\,
            I => \N__22425\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__22431\,
            I => \N__22422\
        );

    \I__2889\ : Odrv12
    port map (
            O => \N__22428\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__22425\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__2887\ : Odrv4
    port map (
            O => \N__22422\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__2886\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__22412\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\
        );

    \I__2884\ : InMux
    port map (
            O => \N__22409\,
            I => \N__22406\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__22406\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\
        );

    \I__2882\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__22400\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\
        );

    \I__2880\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__22394\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__2878\ : InMux
    port map (
            O => \N__22391\,
            I => \N__22388\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__22388\,
            I => \N__22385\
        );

    \I__2876\ : Odrv12
    port map (
            O => \N__22385\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__22382\,
            I => \N__22379\
        );

    \I__2874\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22376\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__22376\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2872\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__22370\,
            I => \N__22367\
        );

    \I__2870\ : Span4Mux_h
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__22364\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__22361\,
            I => \N__22358\
        );

    \I__2867\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__22355\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2865\ : InMux
    port map (
            O => \N__22352\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2864\ : IoInMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__2862\ : Span4Mux_s0_v
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__2861\ : Span4Mux_v
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__2860\ : Sp12to4
    port map (
            O => \N__22337\,
            I => \N__22334\
        );

    \I__2859\ : Span12Mux_h
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__2858\ : Odrv12
    port map (
            O => \N__22331\,
            I => pwm_output_c
        );

    \I__2857\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__2855\ : Odrv12
    port map (
            O => \N__22322\,
            I => il_min_comp1_c
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__22319\,
            I => \N__22315\
        );

    \I__2853\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22312\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22315\,
            I => \N__22309\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__22312\,
            I => \N__22305\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__22309\,
            I => \N__22302\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22308\,
            I => \N__22299\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__22305\,
            I => \N__22294\
        );

    \I__2847\ : Span4Mux_h
    port map (
            O => \N__22302\,
            I => \N__22289\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__22299\,
            I => \N__22289\
        );

    \I__2845\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22284\
        );

    \I__2844\ : InMux
    port map (
            O => \N__22297\,
            I => \N__22284\
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__22294\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__22289\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__22284\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2840\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__22274\,
            I => \N__22271\
        );

    \I__2838\ : Odrv12
    port map (
            O => \N__22271\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22265\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__22265\,
            I => \N__22262\
        );

    \I__2835\ : Odrv12
    port map (
            O => \N__22262\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__22259\,
            I => \N__22256\
        );

    \I__2833\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22253\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__22253\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2831\ : InMux
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__22247\,
            I => \N__22244\
        );

    \I__2829\ : Odrv12
    port map (
            O => \N__22244\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__22241\,
            I => \N__22238\
        );

    \I__2827\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22235\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__22235\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2825\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22229\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__22229\,
            I => \N__22226\
        );

    \I__2823\ : Span4Mux_h
    port map (
            O => \N__22226\,
            I => \N__22223\
        );

    \I__2822\ : Span4Mux_h
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__22220\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__2819\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__22211\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2817\ : InMux
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__2815\ : Span4Mux_h
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__22199\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__2812\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__22190\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2810\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__2808\ : Odrv12
    port map (
            O => \N__22181\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__22172\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__2803\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__2801\ : Odrv4
    port map (
            O => \N__22160\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__2800\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22154\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__22154\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22148\,
            I => \N__22145\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__2795\ : Odrv12
    port map (
            O => \N__22142\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__2794\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22136\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__22136\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__22133\,
            I => \elapsed_time_ns_1_RNI40CED1_0_17_cascade_\
        );

    \I__2791\ : InMux
    port map (
            O => \N__22130\,
            I => \N__22127\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__22127\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__22124\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__22121\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_\
        );

    \I__2787\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22115\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__22115\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24\
        );

    \I__2785\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22109\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__22109\,
            I => \N__22106\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__22106\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__22103\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__2779\ : Odrv12
    port map (
            O => \N__22094\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__22091\,
            I => \N__22088\
        );

    \I__2777\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22085\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__22082\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2774\ : InMux
    port map (
            O => \N__22079\,
            I => \N__22076\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__22076\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__2770\ : Span4Mux_h
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__22064\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__22058\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__22055\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__22052\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16_cascade_\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__22049\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_\
        );

    \I__2763\ : InMux
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__22043\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2\
        );

    \I__2761\ : InMux
    port map (
            O => \N__22040\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\
        );

    \I__2760\ : InMux
    port map (
            O => \N__22037\,
            I => \bfn_8_18_0_\
        );

    \I__2759\ : InMux
    port map (
            O => \N__22034\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\
        );

    \I__2758\ : InMux
    port map (
            O => \N__22031\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\
        );

    \I__2757\ : InMux
    port map (
            O => \N__22028\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\
        );

    \I__2756\ : InMux
    port map (
            O => \N__22025\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\
        );

    \I__2755\ : InMux
    port map (
            O => \N__22022\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\
        );

    \I__2754\ : InMux
    port map (
            O => \N__22019\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\
        );

    \I__2753\ : InMux
    port map (
            O => \N__22016\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_31\
        );

    \I__2752\ : InMux
    port map (
            O => \N__22013\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\
        );

    \I__2751\ : InMux
    port map (
            O => \N__22010\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22007\,
            I => \bfn_8_17_0_\
        );

    \I__2749\ : InMux
    port map (
            O => \N__22004\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\
        );

    \I__2748\ : InMux
    port map (
            O => \N__22001\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\
        );

    \I__2747\ : InMux
    port map (
            O => \N__21998\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\
        );

    \I__2746\ : InMux
    port map (
            O => \N__21995\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\
        );

    \I__2745\ : InMux
    port map (
            O => \N__21992\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\
        );

    \I__2744\ : InMux
    port map (
            O => \N__21989\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\
        );

    \I__2743\ : InMux
    port map (
            O => \N__21986\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\
        );

    \I__2742\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21980\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21977\
        );

    \I__2740\ : Odrv4
    port map (
            O => \N__21977\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\
        );

    \I__2739\ : InMux
    port map (
            O => \N__21974\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\
        );

    \I__2738\ : InMux
    port map (
            O => \N__21971\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\
        );

    \I__2737\ : InMux
    port map (
            O => \N__21968\,
            I => \N__21965\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__21965\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\
        );

    \I__2735\ : InMux
    port map (
            O => \N__21962\,
            I => \bfn_8_16_0_\
        );

    \I__2734\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__21956\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\
        );

    \I__2732\ : InMux
    port map (
            O => \N__21953\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\
        );

    \I__2731\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__21947\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\
        );

    \I__2729\ : InMux
    port map (
            O => \N__21944\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\
        );

    \I__2728\ : InMux
    port map (
            O => \N__21941\,
            I => \N__21938\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__21935\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\
        );

    \I__2725\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__2723\ : Odrv4
    port map (
            O => \N__21926\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_11\
        );

    \I__2722\ : InMux
    port map (
            O => \N__21923\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\
        );

    \I__2721\ : InMux
    port map (
            O => \N__21920\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\
        );

    \I__2720\ : InMux
    port map (
            O => \N__21917\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\
        );

    \I__2719\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21910\
        );

    \I__2718\ : InMux
    port map (
            O => \N__21913\,
            I => \N__21907\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__21910\,
            I => \N__21904\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__21907\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__2715\ : Odrv4
    port map (
            O => \N__21904\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__2714\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21896\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__21896\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\
        );

    \I__2712\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__21890\,
            I => \N__21886\
        );

    \I__2710\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21883\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__21886\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__21883\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__2707\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__21875\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\
        );

    \I__2705\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21869\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__21869\,
            I => \N__21865\
        );

    \I__2703\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21862\
        );

    \I__2702\ : Odrv12
    port map (
            O => \N__21865\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__21862\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__2700\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__21854\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\
        );

    \I__2698\ : InMux
    port map (
            O => \N__21851\,
            I => \N__21848\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__21848\,
            I => \N__21845\
        );

    \I__2696\ : Span4Mux_v
    port map (
            O => \N__21845\,
            I => \N__21841\
        );

    \I__2695\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21838\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__21841\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__21838\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__2692\ : InMux
    port map (
            O => \N__21833\,
            I => \N__21830\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__21830\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\
        );

    \I__2690\ : InMux
    port map (
            O => \N__21827\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\
        );

    \I__2689\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21821\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__21821\,
            I => \N__21818\
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__21818\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__2686\ : InMux
    port map (
            O => \N__21815\,
            I => \N__21810\
        );

    \I__2685\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21807\
        );

    \I__2684\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21804\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__21810\,
            I => \N__21799\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__21807\,
            I => \N__21799\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__21804\,
            I => \N__21794\
        );

    \I__2680\ : Span4Mux_v
    port map (
            O => \N__21799\,
            I => \N__21794\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__21794\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__2678\ : InMux
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__2676\ : Odrv4
    port map (
            O => \N__21785\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__21782\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_\
        );

    \I__2674\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__21776\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__21773\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_\
        );

    \I__2671\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__21767\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__2669\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__21761\,
            I => \current_shift_inst.PI_CTRL.N_62\
        );

    \I__2667\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__21755\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\
        );

    \I__2665\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__21749\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__21746\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_\
        );

    \I__2662\ : IoInMux
    port map (
            O => \N__21743\,
            I => \N__21740\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__2660\ : IoSpan4Mux
    port map (
            O => \N__21737\,
            I => \N__21734\
        );

    \I__2659\ : Span4Mux_s2_v
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__21731\,
            I => \delay_measurement_inst.delay_hc_timer.N_432_i\
        );

    \I__2657\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21725\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__2655\ : Odrv12
    port map (
            O => \N__21722\,
            I => il_max_comp1_c
        );

    \I__2654\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21713\
        );

    \I__2652\ : Span4Mux_h
    port map (
            O => \N__21713\,
            I => \N__21710\
        );

    \I__2651\ : Span4Mux_v
    port map (
            O => \N__21710\,
            I => \N__21707\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__21707\,
            I => il_max_comp2_c
        );

    \I__2649\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__2647\ : Span12Mux_h
    port map (
            O => \N__21698\,
            I => \N__21695\
        );

    \I__2646\ : Odrv12
    port map (
            O => \N__21695\,
            I => il_min_comp2_c
        );

    \I__2645\ : InMux
    port map (
            O => \N__21692\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__2644\ : InMux
    port map (
            O => \N__21689\,
            I => \bfn_7_16_0_\
        );

    \I__2643\ : InMux
    port map (
            O => \N__21686\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__2642\ : InMux
    port map (
            O => \N__21683\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__2641\ : InMux
    port map (
            O => \N__21680\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__2640\ : InMux
    port map (
            O => \N__21677\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__2639\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__21671\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__2637\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__2635\ : Odrv12
    port map (
            O => \N__21662\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__2634\ : InMux
    port map (
            O => \N__21659\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__2633\ : InMux
    port map (
            O => \N__21656\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__2632\ : InMux
    port map (
            O => \N__21653\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__2631\ : InMux
    port map (
            O => \N__21650\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__2630\ : InMux
    port map (
            O => \N__21647\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__2629\ : InMux
    port map (
            O => \N__21644\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__2628\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21638\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__21638\,
            I => \current_shift_inst.PI_CTRL.N_74_16\
        );

    \I__2626\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21629\
        );

    \I__2625\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21629\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__21629\,
            I => \current_shift_inst.PI_CTRL.N_74_21\
        );

    \I__2623\ : InMux
    port map (
            O => \N__21626\,
            I => \N__21620\
        );

    \I__2622\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21620\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__21620\,
            I => \current_shift_inst.PI_CTRL.N_72\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__21617\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1_cascade_\
        );

    \I__2619\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__21611\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__21608\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_\
        );

    \I__2616\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21602\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__21602\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__21599\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__21596\,
            I => \current_shift_inst.PI_CTRL.N_74_16_cascade_\
        );

    \I__2612\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21590\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__21590\,
            I => \N__21587\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__21587\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2609\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21581\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__21581\,
            I => \N__21578\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__21578\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2606\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21572\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__21572\,
            I => \N__21569\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__21569\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2603\ : InMux
    port map (
            O => \N__21566\,
            I => \N__21563\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__21563\,
            I => \N__21560\
        );

    \I__2601\ : Odrv4
    port map (
            O => \N__21560\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2600\ : InMux
    port map (
            O => \N__21557\,
            I => \N__21554\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__21554\,
            I => \N__21551\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__21551\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2597\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21545\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__21545\,
            I => \N__21542\
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__21542\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2594\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21536\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__21536\,
            I => \N__21533\
        );

    \I__2592\ : Span4Mux_h
    port map (
            O => \N__21533\,
            I => \N__21530\
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__21530\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__21527\,
            I => \N__21516\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__21526\,
            I => \N__21512\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__21525\,
            I => \N__21508\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__21524\,
            I => \N__21504\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__21523\,
            I => \N__21500\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__21522\,
            I => \N__21496\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__21521\,
            I => \N__21492\
        );

    \I__2583\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21472\
        );

    \I__2582\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21472\
        );

    \I__2581\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21472\
        );

    \I__2580\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21472\
        );

    \I__2579\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21472\
        );

    \I__2578\ : InMux
    port map (
            O => \N__21511\,
            I => \N__21472\
        );

    \I__2577\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21472\
        );

    \I__2576\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21472\
        );

    \I__2575\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21455\
        );

    \I__2574\ : InMux
    port map (
            O => \N__21503\,
            I => \N__21455\
        );

    \I__2573\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21455\
        );

    \I__2572\ : InMux
    port map (
            O => \N__21499\,
            I => \N__21455\
        );

    \I__2571\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21455\
        );

    \I__2570\ : InMux
    port map (
            O => \N__21495\,
            I => \N__21455\
        );

    \I__2569\ : InMux
    port map (
            O => \N__21492\,
            I => \N__21455\
        );

    \I__2568\ : InMux
    port map (
            O => \N__21491\,
            I => \N__21455\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__21490\,
            I => \N__21452\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__21489\,
            I => \N__21448\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__21472\,
            I => \N__21442\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__21455\,
            I => \N__21442\
        );

    \I__2563\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21433\
        );

    \I__2562\ : InMux
    port map (
            O => \N__21451\,
            I => \N__21433\
        );

    \I__2561\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21433\
        );

    \I__2560\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21433\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__21442\,
            I => \N__21428\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__21433\,
            I => \N__21428\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__21428\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__2556\ : InMux
    port map (
            O => \N__21425\,
            I => \N__21422\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__21422\,
            I => \N__21419\
        );

    \I__2554\ : Odrv12
    port map (
            O => \N__21419\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2553\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21413\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__21413\,
            I => \N__21410\
        );

    \I__2551\ : Odrv12
    port map (
            O => \N__21410\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__2550\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21404\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__2548\ : Odrv12
    port map (
            O => \N__21401\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__21398\,
            I => \N__21395\
        );

    \I__2546\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21392\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21389\
        );

    \I__2544\ : Odrv12
    port map (
            O => \N__21389\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__2543\ : ClkMux
    port map (
            O => \N__21386\,
            I => \N__21380\
        );

    \I__2542\ : ClkMux
    port map (
            O => \N__21385\,
            I => \N__21380\
        );

    \I__2541\ : GlobalMux
    port map (
            O => \N__21380\,
            I => \N__21377\
        );

    \I__2540\ : gio2CtrlBuf
    port map (
            O => \N__21377\,
            I => delay_hc_input_c_g
        );

    \I__2539\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21371\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__2537\ : Glb2LocalMux
    port map (
            O => \N__21368\,
            I => \N__21365\
        );

    \I__2536\ : GlobalMux
    port map (
            O => \N__21365\,
            I => clk_12mhz
        );

    \I__2535\ : IoInMux
    port map (
            O => \N__21362\,
            I => \N__21359\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__21359\,
            I => \N__21356\
        );

    \I__2533\ : IoSpan4Mux
    port map (
            O => \N__21356\,
            I => \N__21353\
        );

    \I__2532\ : Span4Mux_s0_v
    port map (
            O => \N__21353\,
            I => \N__21350\
        );

    \I__2531\ : Odrv4
    port map (
            O => \N__21350\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2530\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21344\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__21344\,
            I => \N__21341\
        );

    \I__2528\ : Span4Mux_h
    port map (
            O => \N__21341\,
            I => \N__21338\
        );

    \I__2527\ : Odrv4
    port map (
            O => \N__21338\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__2526\ : InMux
    port map (
            O => \N__21335\,
            I => \N__21332\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N__21329\
        );

    \I__2524\ : Span4Mux_h
    port map (
            O => \N__21329\,
            I => \N__21326\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__21326\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__2522\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21320\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__21320\,
            I => \N__21317\
        );

    \I__2520\ : Odrv12
    port map (
            O => \N__21317\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__21314\,
            I => \N__21310\
        );

    \I__2518\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21307\
        );

    \I__2517\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21304\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__21307\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__21304\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2514\ : InMux
    port map (
            O => \N__21299\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2513\ : InMux
    port map (
            O => \N__21296\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21287\
        );

    \I__2511\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21287\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__21287\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2509\ : InMux
    port map (
            O => \N__21284\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21281\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2507\ : InMux
    port map (
            O => \N__21278\,
            I => \N__21274\
        );

    \I__2506\ : InMux
    port map (
            O => \N__21277\,
            I => \N__21266\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__21274\,
            I => \N__21261\
        );

    \I__2504\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21254\
        );

    \I__2503\ : InMux
    port map (
            O => \N__21272\,
            I => \N__21254\
        );

    \I__2502\ : InMux
    port map (
            O => \N__21271\,
            I => \N__21254\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21270\,
            I => \N__21248\
        );

    \I__2500\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21248\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__21266\,
            I => \N__21245\
        );

    \I__2498\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21240\
        );

    \I__2497\ : InMux
    port map (
            O => \N__21264\,
            I => \N__21240\
        );

    \I__2496\ : Span4Mux_h
    port map (
            O => \N__21261\,
            I => \N__21237\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__21254\,
            I => \N__21234\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21231\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__21248\,
            I => \N__21226\
        );

    \I__2492\ : Span4Mux_h
    port map (
            O => \N__21245\,
            I => \N__21226\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__21240\,
            I => \N__21223\
        );

    \I__2490\ : Span4Mux_v
    port map (
            O => \N__21237\,
            I => \N__21216\
        );

    \I__2489\ : Span4Mux_h
    port map (
            O => \N__21234\,
            I => \N__21216\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__21231\,
            I => \N__21216\
        );

    \I__2487\ : Span4Mux_v
    port map (
            O => \N__21226\,
            I => \N__21213\
        );

    \I__2486\ : Odrv12
    port map (
            O => \N__21223\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2485\ : Odrv4
    port map (
            O => \N__21216\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__21213\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21203\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__21203\,
            I => \N__21199\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21196\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__21199\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21196\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2478\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__21188\,
            I => \N__21184\
        );

    \I__2476\ : InMux
    port map (
            O => \N__21187\,
            I => \N__21181\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__21184\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__21181\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__21176\,
            I => \N__21173\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21170\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21170\,
            I => \N__21166\
        );

    \I__2470\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21163\
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__21166\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__21163\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__21158\,
            I => \N__21154\
        );

    \I__2466\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21151\
        );

    \I__2465\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21148\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__21151\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__21148\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2462\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21140\,
            I => \N__21136\
        );

    \I__2460\ : InMux
    port map (
            O => \N__21139\,
            I => \N__21133\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__21136\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__21133\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__21128\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\
        );

    \I__2456\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21122\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__21122\,
            I => \N__21118\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21121\,
            I => \N__21115\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__21118\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__21115\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2451\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21107\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__21107\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__2448\ : InMux
    port map (
            O => \N__21101\,
            I => \N__21097\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21094\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__21097\,
            I => \N__21089\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__21094\,
            I => \N__21089\
        );

    \I__2444\ : Odrv4
    port map (
            O => \N__21089\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2443\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21083\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__21083\,
            I => \N__21079\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21082\,
            I => \N__21076\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__21079\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__21076\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2438\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21068\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__21068\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__2436\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21059\
        );

    \I__2435\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21059\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__21059\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2433\ : InMux
    port map (
            O => \N__21056\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2432\ : InMux
    port map (
            O => \N__21053\,
            I => \N__21050\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__2430\ : Span4Mux_h
    port map (
            O => \N__21047\,
            I => \N__21043\
        );

    \I__2429\ : InMux
    port map (
            O => \N__21046\,
            I => \N__21040\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__21043\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__21040\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2426\ : InMux
    port map (
            O => \N__21035\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2425\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21029\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__2423\ : Span4Mux_h
    port map (
            O => \N__21026\,
            I => \N__21022\
        );

    \I__2422\ : InMux
    port map (
            O => \N__21025\,
            I => \N__21019\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__21022\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__21019\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2419\ : InMux
    port map (
            O => \N__21014\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2418\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21005\
        );

    \I__2417\ : InMux
    port map (
            O => \N__21010\,
            I => \N__21005\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__21005\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2415\ : InMux
    port map (
            O => \N__21002\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2414\ : InMux
    port map (
            O => \N__20999\,
            I => \N__20993\
        );

    \I__2413\ : InMux
    port map (
            O => \N__20998\,
            I => \N__20993\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__20993\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2411\ : InMux
    port map (
            O => \N__20990\,
            I => \bfn_5_13_0_\
        );

    \I__2410\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20981\
        );

    \I__2409\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20981\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__20981\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2407\ : InMux
    port map (
            O => \N__20978\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2406\ : InMux
    port map (
            O => \N__20975\,
            I => \N__20969\
        );

    \I__2405\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20969\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__20969\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2403\ : InMux
    port map (
            O => \N__20966\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2402\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20957\
        );

    \I__2401\ : InMux
    port map (
            O => \N__20962\,
            I => \N__20957\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__20957\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2399\ : InMux
    port map (
            O => \N__20954\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2398\ : InMux
    port map (
            O => \N__20951\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2397\ : InMux
    port map (
            O => \N__20948\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__20945\,
            I => \N__20942\
        );

    \I__2395\ : InMux
    port map (
            O => \N__20942\,
            I => \N__20939\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__20939\,
            I => \N__20935\
        );

    \I__2393\ : InMux
    port map (
            O => \N__20938\,
            I => \N__20932\
        );

    \I__2392\ : Span4Mux_h
    port map (
            O => \N__20935\,
            I => \N__20929\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__20932\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2390\ : Odrv4
    port map (
            O => \N__20929\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2389\ : InMux
    port map (
            O => \N__20924\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__20921\,
            I => \N__20917\
        );

    \I__2387\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20914\
        );

    \I__2386\ : InMux
    port map (
            O => \N__20917\,
            I => \N__20911\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__20914\,
            I => \N__20908\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__20911\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__20908\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2382\ : InMux
    port map (
            O => \N__20903\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2381\ : InMux
    port map (
            O => \N__20900\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2380\ : InMux
    port map (
            O => \N__20897\,
            I => \bfn_5_12_0_\
        );

    \I__2379\ : InMux
    port map (
            O => \N__20894\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2378\ : InMux
    port map (
            O => \N__20891\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__20888\,
            I => \N__20884\
        );

    \I__2376\ : InMux
    port map (
            O => \N__20887\,
            I => \N__20881\
        );

    \I__2375\ : InMux
    port map (
            O => \N__20884\,
            I => \N__20878\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__20881\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__20878\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2372\ : InMux
    port map (
            O => \N__20873\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2371\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20864\
        );

    \I__2370\ : InMux
    port map (
            O => \N__20869\,
            I => \N__20864\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__20864\,
            I => \N__20860\
        );

    \I__2368\ : InMux
    port map (
            O => \N__20863\,
            I => \N__20857\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__20860\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__20857\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2365\ : InMux
    port map (
            O => \N__20852\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2364\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20845\
        );

    \I__2363\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20842\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__20845\,
            I => \N__20839\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__20842\,
            I => \N__20836\
        );

    \I__2360\ : Span4Mux_h
    port map (
            O => \N__20839\,
            I => \N__20831\
        );

    \I__2359\ : Span4Mux_h
    port map (
            O => \N__20836\,
            I => \N__20828\
        );

    \I__2358\ : InMux
    port map (
            O => \N__20835\,
            I => \N__20823\
        );

    \I__2357\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20823\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__20831\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__20828\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__20823\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2353\ : InMux
    port map (
            O => \N__20816\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__2351\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__20804\,
            I => \N__20799\
        );

    \I__2348\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20796\
        );

    \I__2347\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20793\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__20799\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__20796\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__20793\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2343\ : InMux
    port map (
            O => \N__20786\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__2341\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20775\
        );

    \I__2340\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20772\
        );

    \I__2339\ : InMux
    port map (
            O => \N__20778\,
            I => \N__20769\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__20775\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__20772\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__20769\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2335\ : InMux
    port map (
            O => \N__20762\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2334\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__2332\ : Span4Mux_h
    port map (
            O => \N__20753\,
            I => \N__20748\
        );

    \I__2331\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20745\
        );

    \I__2330\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20742\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__20748\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__20745\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__20742\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2326\ : InMux
    port map (
            O => \N__20735\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__20732\,
            I => \N__20728\
        );

    \I__2324\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20724\
        );

    \I__2323\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20721\
        );

    \I__2322\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20718\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__20724\,
            I => \N__20715\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__20721\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__20718\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__20715\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2317\ : InMux
    port map (
            O => \N__20708\,
            I => \bfn_5_11_0_\
        );

    \I__2316\ : InMux
    port map (
            O => \N__20705\,
            I => \N__20701\
        );

    \I__2315\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20698\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__20701\,
            I => \N__20692\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__20698\,
            I => \N__20692\
        );

    \I__2312\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20689\
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__20692\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__20689\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2309\ : InMux
    port map (
            O => \N__20684\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2308\ : InMux
    port map (
            O => \N__20681\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2307\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__20675\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__20672\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\
        );

    \I__2304\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20658\
        );

    \I__2303\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20653\
        );

    \I__2302\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20653\
        );

    \I__2301\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20646\
        );

    \I__2300\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20646\
        );

    \I__2299\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20646\
        );

    \I__2298\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20643\
        );

    \I__2297\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20638\
        );

    \I__2296\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20638\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__20658\,
            I => \N__20635\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__20653\,
            I => \N__20632\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__20646\,
            I => \N__20625\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__20643\,
            I => \N__20625\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__20638\,
            I => \N__20625\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__20635\,
            I => \N__20622\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__20632\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__20625\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__20622\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2286\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20612\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__20612\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2284\ : InMux
    port map (
            O => \N__20609\,
            I => \N__20606\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__20606\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2282\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20600\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__20600\,
            I => \N__20597\
        );

    \I__2280\ : Span4Mux_h
    port map (
            O => \N__20597\,
            I => \N__20594\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__20594\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__2278\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20588\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__20588\,
            I => \N__20585\
        );

    \I__2276\ : Span4Mux_h
    port map (
            O => \N__20585\,
            I => \N__20582\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__20582\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__2274\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20576\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__20576\,
            I => \N__20573\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__20573\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2271\ : InMux
    port map (
            O => \N__20570\,
            I => \N__20567\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__20567\,
            I => \N__20564\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__20564\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2268\ : InMux
    port map (
            O => \N__20561\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__2267\ : InMux
    port map (
            O => \N__20558\,
            I => \N__20555\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__20555\,
            I => \N__20552\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__20552\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2264\ : InMux
    port map (
            O => \N__20549\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2263\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20543\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__20543\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__20540\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\
        );

    \I__2260\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20534\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__20534\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__20531\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\
        );

    \I__2257\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20525\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__20525\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__20522\,
            I => \N__20517\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__20521\,
            I => \N__20512\
        );

    \I__2253\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20507\
        );

    \I__2252\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20507\
        );

    \I__2251\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20499\
        );

    \I__2250\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20499\
        );

    \I__2249\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20499\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__20507\,
            I => \N__20496\
        );

    \I__2247\ : InMux
    port map (
            O => \N__20506\,
            I => \N__20492\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__20499\,
            I => \N__20487\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__20496\,
            I => \N__20487\
        );

    \I__2244\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20484\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__20492\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__20487\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__20484\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2240\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20474\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__20474\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__20471\,
            I => \N__20468\
        );

    \I__2237\ : InMux
    port map (
            O => \N__20468\,
            I => \N__20465\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__20465\,
            I => \N__20462\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__20462\,
            I => \N__20459\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__20459\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9\
        );

    \I__2233\ : InMux
    port map (
            O => \N__20456\,
            I => \N__20453\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__20453\,
            I => \N__20448\
        );

    \I__2231\ : InMux
    port map (
            O => \N__20452\,
            I => \N__20445\
        );

    \I__2230\ : InMux
    port map (
            O => \N__20451\,
            I => \N__20442\
        );

    \I__2229\ : Span4Mux_h
    port map (
            O => \N__20448\,
            I => \N__20439\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__20445\,
            I => pwm_duty_input_9
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__20442\,
            I => pwm_duty_input_9
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__20439\,
            I => pwm_duty_input_9
        );

    \I__2225\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20429\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__20429\,
            I => \N__20425\
        );

    \I__2223\ : InMux
    port map (
            O => \N__20428\,
            I => \N__20422\
        );

    \I__2222\ : Span4Mux_v
    port map (
            O => \N__20425\,
            I => \N__20417\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__20422\,
            I => \N__20417\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__20417\,
            I => \N__20413\
        );

    \I__2219\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20410\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__20413\,
            I => pwm_duty_input_7
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__20410\,
            I => pwm_duty_input_7
        );

    \I__2216\ : InMux
    port map (
            O => \N__20405\,
            I => \N__20401\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__20404\,
            I => \N__20398\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__20401\,
            I => \N__20394\
        );

    \I__2213\ : InMux
    port map (
            O => \N__20398\,
            I => \N__20391\
        );

    \I__2212\ : InMux
    port map (
            O => \N__20397\,
            I => \N__20388\
        );

    \I__2211\ : Span4Mux_h
    port map (
            O => \N__20394\,
            I => \N__20385\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__20391\,
            I => pwm_duty_input_6
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__20388\,
            I => pwm_duty_input_6
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__20385\,
            I => pwm_duty_input_6
        );

    \I__2207\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__20375\,
            I => \N__20370\
        );

    \I__2205\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20367\
        );

    \I__2204\ : InMux
    port map (
            O => \N__20373\,
            I => \N__20364\
        );

    \I__2203\ : Span4Mux_v
    port map (
            O => \N__20370\,
            I => \N__20361\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__20367\,
            I => pwm_duty_input_8
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__20364\,
            I => pwm_duty_input_8
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__20361\,
            I => pwm_duty_input_8
        );

    \I__2199\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__20351\,
            I => \N__20346\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20343\
        );

    \I__2196\ : InMux
    port map (
            O => \N__20349\,
            I => \N__20340\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__20346\,
            I => \N__20337\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__20343\,
            I => pwm_duty_input_3
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__20340\,
            I => pwm_duty_input_3
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__20337\,
            I => pwm_duty_input_3
        );

    \I__2191\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20325\
        );

    \I__2190\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20322\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20328\,
            I => \N__20319\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__20325\,
            I => \N__20316\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__20322\,
            I => \N__20313\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__20319\,
            I => \N__20310\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__20316\,
            I => pwm_duty_input_4
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__20313\,
            I => pwm_duty_input_4
        );

    \I__2183\ : Odrv12
    port map (
            O => \N__20310\,
            I => pwm_duty_input_4
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__20303\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20297\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__20297\,
            I => \N__20293\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20290\
        );

    \I__2178\ : Span4Mux_v
    port map (
            O => \N__20293\,
            I => \N__20285\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__20290\,
            I => \N__20285\
        );

    \I__2176\ : Span4Mux_h
    port map (
            O => \N__20285\,
            I => \N__20281\
        );

    \I__2175\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20278\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__20281\,
            I => pwm_duty_input_5
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__20278\,
            I => pwm_duty_input_5
        );

    \I__2172\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20251\
        );

    \I__2171\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20251\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20251\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20251\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20251\
        );

    \I__2167\ : InMux
    port map (
            O => \N__20268\,
            I => \N__20251\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20242\
        );

    \I__2165\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20242\
        );

    \I__2164\ : InMux
    port map (
            O => \N__20265\,
            I => \N__20242\
        );

    \I__2163\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20242\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__20251\,
            I => \N__20237\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__20242\,
            I => \N__20237\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__20237\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__20234\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__2157\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20224\
        );

    \I__2156\ : InMux
    port map (
            O => \N__20227\,
            I => \N__20221\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__20224\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__20221\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__20216\,
            I => \N__20213\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20213\,
            I => \N__20210\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__20210\,
            I => \current_shift_inst.PI_CTRL.N_155\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__20207\,
            I => \N__20203\
        );

    \I__2149\ : InMux
    port map (
            O => \N__20206\,
            I => \N__20200\
        );

    \I__2148\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20197\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__20200\,
            I => \N__20191\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__20197\,
            I => \N__20191\
        );

    \I__2145\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20188\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__20191\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__20188\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20180\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__20180\,
            I => \current_shift_inst.PI_CTRL.N_149\
        );

    \I__2140\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__20174\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__2138\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20168\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__20168\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__20165\,
            I => \N__20162\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20159\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__20159\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__20156\,
            I => \N__20153\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20153\,
            I => \N__20150\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__20150\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__2130\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20144\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__20144\,
            I => \N__20141\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__20141\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__2127\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20135\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__20135\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__2125\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20129\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__20129\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__2123\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20104\
        );

    \I__2122\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20104\
        );

    \I__2121\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20104\
        );

    \I__2120\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20104\
        );

    \I__2119\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20104\
        );

    \I__2118\ : InMux
    port map (
            O => \N__20121\,
            I => \N__20104\
        );

    \I__2117\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20095\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20095\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20095\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20117\,
            I => \N__20095\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__20092\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__20095\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__20092\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__20087\,
            I => \N__20084\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__20081\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__20078\,
            I => \N__20070\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__20077\,
            I => \N__20059\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__20076\,
            I => \N__20056\
        );

    \I__2104\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20047\
        );

    \I__2103\ : InMux
    port map (
            O => \N__20074\,
            I => \N__20047\
        );

    \I__2102\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20047\
        );

    \I__2101\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20047\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__20069\,
            I => \N__20042\
        );

    \I__2099\ : InMux
    port map (
            O => \N__20068\,
            I => \N__20035\
        );

    \I__2098\ : InMux
    port map (
            O => \N__20067\,
            I => \N__20035\
        );

    \I__2097\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20035\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20022\
        );

    \I__2095\ : InMux
    port map (
            O => \N__20064\,
            I => \N__20022\
        );

    \I__2094\ : InMux
    port map (
            O => \N__20063\,
            I => \N__20022\
        );

    \I__2093\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20022\
        );

    \I__2092\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20022\
        );

    \I__2091\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20022\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__20047\,
            I => \N__20019\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20046\,
            I => \N__20014\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20045\,
            I => \N__20014\
        );

    \I__2087\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20011\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__20035\,
            I => \N__20008\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__20022\,
            I => \N__20005\
        );

    \I__2084\ : Span4Mux_h
    port map (
            O => \N__20019\,
            I => \N__19984\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__19984\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__20011\,
            I => \N__19979\
        );

    \I__2081\ : Span4Mux_s1_h
    port map (
            O => \N__20008\,
            I => \N__19979\
        );

    \I__2080\ : Span4Mux_h
    port map (
            O => \N__20005\,
            I => \N__19976\
        );

    \I__2079\ : InMux
    port map (
            O => \N__20004\,
            I => \N__19973\
        );

    \I__2078\ : InMux
    port map (
            O => \N__20003\,
            I => \N__19956\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20002\,
            I => \N__19956\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19956\
        );

    \I__2075\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19956\
        );

    \I__2074\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19956\
        );

    \I__2073\ : InMux
    port map (
            O => \N__19998\,
            I => \N__19956\
        );

    \I__2072\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19956\
        );

    \I__2071\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19956\
        );

    \I__2070\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19941\
        );

    \I__2069\ : InMux
    port map (
            O => \N__19994\,
            I => \N__19941\
        );

    \I__2068\ : InMux
    port map (
            O => \N__19993\,
            I => \N__19941\
        );

    \I__2067\ : InMux
    port map (
            O => \N__19992\,
            I => \N__19941\
        );

    \I__2066\ : InMux
    port map (
            O => \N__19991\,
            I => \N__19941\
        );

    \I__2065\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19941\
        );

    \I__2064\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19941\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__19984\,
            I => \N__19936\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__19979\,
            I => \N__19936\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__19976\,
            I => \N_19_1\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__19973\,
            I => \N_19_1\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__19956\,
            I => \N_19_1\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__19941\,
            I => \N_19_1\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__19936\,
            I => \N_19_1\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__19925\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__2055\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19916\
        );

    \I__2054\ : InMux
    port map (
            O => \N__19921\,
            I => \N__19916\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__19916\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__2052\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19910\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__19910\,
            I => \N__19906\
        );

    \I__2050\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19903\
        );

    \I__2049\ : Span4Mux_s3_h
    port map (
            O => \N__19906\,
            I => \N__19900\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__19903\,
            I => pwm_duty_input_2
        );

    \I__2047\ : Odrv4
    port map (
            O => \N__19900\,
            I => pwm_duty_input_2
        );

    \I__2046\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19889\
        );

    \I__2045\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19889\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__19889\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__2043\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__19883\,
            I => \N__19879\
        );

    \I__2041\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19876\
        );

    \I__2040\ : Span4Mux_s3_h
    port map (
            O => \N__19879\,
            I => \N__19873\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__19876\,
            I => pwm_duty_input_1
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__19873\,
            I => pwm_duty_input_1
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__19868\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__2036\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__19862\,
            I => \N__19859\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__19859\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__19856\,
            I => \N__19850\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__19855\,
            I => \N__19846\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__19854\,
            I => \N__19843\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__19853\,
            I => \N__19840\
        );

    \I__2029\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19835\
        );

    \I__2028\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19835\
        );

    \I__2027\ : InMux
    port map (
            O => \N__19846\,
            I => \N__19828\
        );

    \I__2026\ : InMux
    port map (
            O => \N__19843\,
            I => \N__19828\
        );

    \I__2025\ : InMux
    port map (
            O => \N__19840\,
            I => \N__19828\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__19835\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__19828\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__2022\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19814\
        );

    \I__2021\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19814\
        );

    \I__2020\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19814\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__19814\,
            I => \current_shift_inst.PI_CTRL.N_154\
        );

    \I__2018\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__19808\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__2016\ : InMux
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__19802\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__2014\ : InMux
    port map (
            O => \N__19799\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__2013\ : InMux
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__19793\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__2011\ : InMux
    port map (
            O => \N__19790\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__2010\ : InMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__19784\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__2008\ : InMux
    port map (
            O => \N__19781\,
            I => \bfn_3_9_0_\
        );

    \I__2007\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19775\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__19772\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__2004\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__19763\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__19760\,
            I => \N__19755\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__19759\,
            I => \N__19750\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__19758\,
            I => \N__19745\
        );

    \I__1998\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19741\
        );

    \I__1997\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19738\
        );

    \I__1996\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19735\
        );

    \I__1995\ : InMux
    port map (
            O => \N__19750\,
            I => \N__19732\
        );

    \I__1994\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19727\
        );

    \I__1993\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19727\
        );

    \I__1992\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19723\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__19744\,
            I => \N__19720\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__19741\,
            I => \N__19714\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__19738\,
            I => \N__19711\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__19735\,
            I => \N__19704\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__19732\,
            I => \N__19704\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__19727\,
            I => \N__19704\
        );

    \I__1985\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19701\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__19723\,
            I => \N__19698\
        );

    \I__1983\ : InMux
    port map (
            O => \N__19720\,
            I => \N__19689\
        );

    \I__1982\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19689\
        );

    \I__1981\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19689\
        );

    \I__1980\ : InMux
    port map (
            O => \N__19717\,
            I => \N__19689\
        );

    \I__1979\ : Span4Mux_h
    port map (
            O => \N__19714\,
            I => \N__19680\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__19711\,
            I => \N__19680\
        );

    \I__1977\ : Span4Mux_h
    port map (
            O => \N__19704\,
            I => \N__19680\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__19701\,
            I => \N__19680\
        );

    \I__1975\ : Span4Mux_h
    port map (
            O => \N__19698\,
            I => \N__19677\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__19689\,
            I => \N__19672\
        );

    \I__1973\ : Span4Mux_s2_h
    port map (
            O => \N__19680\,
            I => \N__19672\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__19677\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__19672\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__1970\ : InMux
    port map (
            O => \N__19667\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__19664\,
            I => \pwm_generator_inst.un1_duty_inputlt3_cascade_\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__19661\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_\
        );

    \I__1967\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__19655\,
            I => \N__19651\
        );

    \I__1965\ : InMux
    port map (
            O => \N__19654\,
            I => \N__19648\
        );

    \I__1964\ : Span4Mux_v
    port map (
            O => \N__19651\,
            I => \N__19645\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__19648\,
            I => pwm_duty_input_0
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__19645\,
            I => pwm_duty_input_0
        );

    \I__1961\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__19637\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__1959\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__19631\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__19628\,
            I => \N__19625\
        );

    \I__1956\ : InMux
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__19622\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__1954\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__19613\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__1950\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__19604\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__1948\ : InMux
    port map (
            O => \N__19601\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__1947\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__19595\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__19592\,
            I => \N__19589\
        );

    \I__1944\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__19586\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__1942\ : InMux
    port map (
            O => \N__19583\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__1941\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__19577\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__19574\,
            I => \N__19571\
        );

    \I__1938\ : InMux
    port map (
            O => \N__19571\,
            I => \N__19568\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__19568\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__1936\ : InMux
    port map (
            O => \N__19565\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__1935\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__19559\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__1933\ : InMux
    port map (
            O => \N__19556\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__1932\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19550\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__19550\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__1930\ : InMux
    port map (
            O => \N__19547\,
            I => \N__19544\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__19544\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__1928\ : InMux
    port map (
            O => \N__19541\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__1927\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__19535\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__1925\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19529\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__19529\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__1923\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__19523\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__1921\ : InMux
    port map (
            O => \N__19520\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__1920\ : InMux
    port map (
            O => \N__19517\,
            I => \N__19514\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__19514\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__1918\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__19508\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__1916\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__19502\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__1914\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__19496\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__1912\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__19490\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__1910\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19484\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__19484\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__1908\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__19478\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__1906\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19472\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__19472\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__1904\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19466\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__19466\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__1902\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__19460\,
            I => \N__19457\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__19457\,
            I => \N__19454\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__19454\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__19451\,
            I => \N__19448\
        );

    \I__1897\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19442\
        );

    \I__1896\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19442\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__19442\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1894\ : InMux
    port map (
            O => \N__19439\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__1893\ : InMux
    port map (
            O => \N__19436\,
            I => \N__19433\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__19433\,
            I => \N__19430\
        );

    \I__1891\ : Span4Mux_v
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__19427\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1889\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19418\
        );

    \I__1888\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19418\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__19418\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__1886\ : InMux
    port map (
            O => \N__19415\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__1885\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19409\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__19409\,
            I => \N__19406\
        );

    \I__1883\ : Span4Mux_h
    port map (
            O => \N__19406\,
            I => \N__19403\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__19403\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__19400\,
            I => \N__19397\
        );

    \I__1880\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19393\
        );

    \I__1879\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19390\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__19393\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__19390\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1876\ : InMux
    port map (
            O => \N__19385\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__1875\ : InMux
    port map (
            O => \N__19382\,
            I => \N__19379\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__19379\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__1872\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__19370\,
            I => \N__19366\
        );

    \I__1870\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__19366\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__19363\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1867\ : InMux
    port map (
            O => \N__19358\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__1865\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__19349\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__1863\ : InMux
    port map (
            O => \N__19346\,
            I => \N__19340\
        );

    \I__1862\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19340\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__19340\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1860\ : InMux
    port map (
            O => \N__19337\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__1859\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__19331\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__1857\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19324\
        );

    \I__1856\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19321\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__19324\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__19321\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1853\ : InMux
    port map (
            O => \N__19316\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__1851\ : InMux
    port map (
            O => \N__19310\,
            I => \N__19307\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__19307\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__1849\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__19301\,
            I => \N__19297\
        );

    \I__1847\ : InMux
    port map (
            O => \N__19300\,
            I => \N__19294\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__19297\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__19294\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__1844\ : InMux
    port map (
            O => \N__19289\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__1843\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__19283\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__1841\ : InMux
    port map (
            O => \N__19280\,
            I => \bfn_2_11_0_\
        );

    \I__1840\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__19274\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__1838\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19266\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19270\,
            I => \N__19263\
        );

    \I__1836\ : InMux
    port map (
            O => \N__19269\,
            I => \N__19260\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__19266\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__19263\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__19260\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1832\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19249\
        );

    \I__1831\ : InMux
    port map (
            O => \N__19252\,
            I => \N__19246\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__19249\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__19246\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__1828\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__19238\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__19235\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19232\,
            I => \N__19228\
        );

    \I__1824\ : InMux
    port map (
            O => \N__19231\,
            I => \N__19225\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__19228\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__19225\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__1821\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__19217\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__19214\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\
        );

    \I__1818\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__19208\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__1816\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19198\
        );

    \I__1815\ : InMux
    port map (
            O => \N__19204\,
            I => \N__19198\
        );

    \I__1814\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19195\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__19198\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__19195\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1811\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__19187\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__1809\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19179\
        );

    \I__1808\ : InMux
    port map (
            O => \N__19183\,
            I => \N__19174\
        );

    \I__1807\ : InMux
    port map (
            O => \N__19182\,
            I => \N__19174\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__19179\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__19174\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__1804\ : InMux
    port map (
            O => \N__19169\,
            I => \N__19165\
        );

    \I__1803\ : InMux
    port map (
            O => \N__19168\,
            I => \N__19162\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__19165\,
            I => \N__19159\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__19162\,
            I => \N__19156\
        );

    \I__1800\ : Span4Mux_v
    port map (
            O => \N__19159\,
            I => \N__19153\
        );

    \I__1799\ : Span4Mux_h
    port map (
            O => \N__19156\,
            I => \N__19150\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__19153\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1797\ : Odrv4
    port map (
            O => \N__19150\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1796\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19142\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__19139\,
            I => \N__19135\
        );

    \I__1793\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19132\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__19135\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__19132\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19127\,
            I => \N__19121\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__19126\,
            I => \N__19117\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__19125\,
            I => \N__19113\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__19124\,
            I => \N__19109\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__19121\,
            I => \N__19106\
        );

    \I__1785\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19092\
        );

    \I__1784\ : InMux
    port map (
            O => \N__19117\,
            I => \N__19092\
        );

    \I__1783\ : InMux
    port map (
            O => \N__19116\,
            I => \N__19092\
        );

    \I__1782\ : InMux
    port map (
            O => \N__19113\,
            I => \N__19092\
        );

    \I__1781\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19092\
        );

    \I__1780\ : InMux
    port map (
            O => \N__19109\,
            I => \N__19092\
        );

    \I__1779\ : Span4Mux_v
    port map (
            O => \N__19106\,
            I => \N__19089\
        );

    \I__1778\ : InMux
    port map (
            O => \N__19105\,
            I => \N__19086\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__19092\,
            I => \N__19083\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__19089\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__19086\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__19083\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__19067\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__19061\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19055\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__19055\,
            I => \rgb_drv_RNOZ0\
        );

    \I__1765\ : InMux
    port map (
            O => \N__19052\,
            I => \N__19049\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__19049\,
            I => \N_38_i_i\
        );

    \I__1763\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19039\
        );

    \I__1762\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19039\
        );

    \I__1761\ : InMux
    port map (
            O => \N__19044\,
            I => \N__19036\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__19039\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__19036\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__1758\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__19028\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19025\,
            I => \N__19021\
        );

    \I__1755\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19018\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__19021\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__19018\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1752\ : InMux
    port map (
            O => \N__19013\,
            I => \N__19007\
        );

    \I__1751\ : InMux
    port map (
            O => \N__19012\,
            I => \N__19007\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__19007\,
            I => \N__19004\
        );

    \I__1749\ : Span4Mux_h
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__19001\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1747\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__18995\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__18992\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\
        );

    \I__1744\ : InMux
    port map (
            O => \N__18989\,
            I => \N__18986\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__18986\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__1742\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18978\
        );

    \I__1741\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18975\
        );

    \I__1740\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18972\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__18978\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__18975\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__18972\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1736\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18962\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__18962\,
            I => \N__18959\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__18959\,
            I => \N__18956\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__18956\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__18953\,
            I => \N__18950\
        );

    \I__1731\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18947\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__18944\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__1728\ : InMux
    port map (
            O => \N__18941\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1727\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18935\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__18935\,
            I => \N__18932\
        );

    \I__1725\ : Span4Mux_v
    port map (
            O => \N__18932\,
            I => \N__18929\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__18929\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1723\ : InMux
    port map (
            O => \N__18926\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__18923\,
            I => \N__18920\
        );

    \I__1721\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__1719\ : Span4Mux_v
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__18911\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1717\ : InMux
    port map (
            O => \N__18908\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1716\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__18899\,
            I => \N__18896\
        );

    \I__1713\ : Odrv4
    port map (
            O => \N__18896\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1712\ : InMux
    port map (
            O => \N__18893\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__1710\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__18878\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__1706\ : InMux
    port map (
            O => \N__18875\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__1705\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__1703\ : Span4Mux_v
    port map (
            O => \N__18866\,
            I => \N__18863\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__18863\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__1701\ : InMux
    port map (
            O => \N__18860\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__1699\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__18851\,
            I => \N__18848\
        );

    \I__1697\ : Odrv12
    port map (
            O => \N__18848\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__1696\ : InMux
    port map (
            O => \N__18845\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__1695\ : InMux
    port map (
            O => \N__18842\,
            I => \bfn_1_12_0_\
        );

    \I__1694\ : InMux
    port map (
            O => \N__18839\,
            I => \N__18836\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__18830\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__1689\ : InMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__18818\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1686\ : InMux
    port map (
            O => \N__18815\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1685\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__18803\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__1680\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__18791\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1677\ : InMux
    port map (
            O => \N__18788\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1676\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__1674\ : Span4Mux_v
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__18776\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__1671\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18767\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__18767\,
            I => \N__18764\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__18764\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1668\ : InMux
    port map (
            O => \N__18761\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1667\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__18755\,
            I => \N__18752\
        );

    \I__1665\ : Span4Mux_v
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__18749\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__1662\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18740\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__1660\ : Span4Mux_v
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__18734\,
            I => \N__18731\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__18731\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1657\ : InMux
    port map (
            O => \N__18728\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1656\ : InMux
    port map (
            O => \N__18725\,
            I => \N__18722\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__18722\,
            I => \N__18719\
        );

    \I__1654\ : Span4Mux_v
    port map (
            O => \N__18719\,
            I => \N__18716\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__18716\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__18713\,
            I => \N__18710\
        );

    \I__1651\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__18707\,
            I => \N__18704\
        );

    \I__1649\ : Span4Mux_h
    port map (
            O => \N__18704\,
            I => \N__18701\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__18701\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__1647\ : InMux
    port map (
            O => \N__18698\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__1646\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__18689\,
            I => \N__18686\
        );

    \I__1643\ : Odrv4
    port map (
            O => \N__18686\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__18683\,
            I => \N__18680\
        );

    \I__1641\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18677\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__18677\,
            I => \N__18674\
        );

    \I__1639\ : Span4Mux_h
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__18671\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__1637\ : InMux
    port map (
            O => \N__18668\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__1636\ : InMux
    port map (
            O => \N__18665\,
            I => \N__18662\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__18662\,
            I => \N__18659\
        );

    \I__1634\ : Span4Mux_v
    port map (
            O => \N__18659\,
            I => \N__18656\
        );

    \I__1633\ : Odrv4
    port map (
            O => \N__18656\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__18653\,
            I => \N__18650\
        );

    \I__1631\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18647\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__18647\,
            I => \N__18644\
        );

    \I__1629\ : Span4Mux_h
    port map (
            O => \N__18644\,
            I => \N__18641\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__18641\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__1627\ : InMux
    port map (
            O => \N__18638\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__1626\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18632\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__18632\,
            I => \N__18629\
        );

    \I__1624\ : Span4Mux_v
    port map (
            O => \N__18629\,
            I => \N__18626\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__18626\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__18623\,
            I => \N__18620\
        );

    \I__1621\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__18617\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__1619\ : InMux
    port map (
            O => \N__18614\,
            I => \bfn_1_11_0_\
        );

    \I__1618\ : InMux
    port map (
            O => \N__18611\,
            I => \bfn_1_9_0_\
        );

    \I__1617\ : InMux
    port map (
            O => \N__18608\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__1616\ : InMux
    port map (
            O => \N__18605\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__1615\ : InMux
    port map (
            O => \N__18602\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__1614\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__1612\ : Span4Mux_v
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__18590\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__18587\,
            I => \N__18584\
        );

    \I__1609\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__18581\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1607\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18575\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__1605\ : Span4Mux_h
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__18569\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1603\ : InMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__18563\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \I__1601\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__18554\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1598\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__18548\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__1596\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__18539\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1593\ : InMux
    port map (
            O => \N__18536\,
            I => \N__18533\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__18533\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__1591\ : InMux
    port map (
            O => \N__18530\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__1590\ : InMux
    port map (
            O => \N__18527\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__1589\ : InMux
    port map (
            O => \N__18524\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__1588\ : InMux
    port map (
            O => \N__18521\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__1587\ : InMux
    port map (
            O => \N__18518\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__1586\ : InMux
    port map (
            O => \N__18515\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__1585\ : InMux
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__1583\ : Odrv4
    port map (
            O => \N__18506\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1582\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__18500\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__1580\ : InMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__18491\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1577\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__18485\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__1575\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__1573\ : Odrv4
    port map (
            O => \N__18476\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1572\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__18470\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__1570\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__18464\,
            I => \N__18461\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__18461\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1567\ : InMux
    port map (
            O => \N__18458\,
            I => \N__18455\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__18455\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__1565\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18449\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__18446\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1562\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__18440\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__1560\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__18431\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1557\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__18425\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__1555\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__1553\ : Span4Mux_h
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__18413\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1551\ : InMux
    port map (
            O => \N__18410\,
            I => \N__18407\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__18407\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__1549\ : IoInMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__1547\ : Span4Mux_s3_v
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__1546\ : Span4Mux_h
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__1545\ : Sp12to4
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__1544\ : Span12Mux_s9_v
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__1543\ : Span12Mux_v
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__1542\ : Odrv12
    port map (
            O => \N__18383\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1541\ : IoInMux
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__1539\ : IoSpan4Mux
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__1538\ : IoSpan4Mux
    port map (
            O => \N__18371\,
            I => \N__18368\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__18368\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_10_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_10_25_0_\
        );

    \IN_MUX_bfv_10_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_10_26_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_3_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_8_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_8\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_16\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_8\,
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_16\,
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_8\,
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_16\,
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_8\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_16\,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_15_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_5_0_\
        );

    \IN_MUX_bfv_15_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_15_6_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_12_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_12_23_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_16_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_16_25_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_7\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_7_16_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18404\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18380\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32402\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_166_i_g\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__33677\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_434_i_g\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21743\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_432_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__37811\,
            CLKHFEN => \N__37813\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__37812\,
            RGB2PWM => \N__19052\,
            RGB1 => rgb_g_wire,
            CURREN => \N__37879\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__19058\,
            RGB0PWM => \N__45728\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21278\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46118\,
            ce => 'H',
            sr => \N__45590\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__19127\,
            in1 => \N__19138\,
            in2 => \_gnd_net_\,
            in3 => \N__20004\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18503\,
            in2 => \_gnd_net_\,
            in3 => \N__18512\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18497\,
            in1 => \N__18488\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18473\,
            in2 => \_gnd_net_\,
            in3 => \N__18482\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18458\,
            in2 => \_gnd_net_\,
            in3 => \N__18467\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18452\,
            in1 => \N__18443\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18428\,
            in2 => \_gnd_net_\,
            in3 => \N__18437\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18410\,
            in2 => \_gnd_net_\,
            in3 => \N__18422\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18566\,
            in2 => \_gnd_net_\,
            in3 => \N__18578\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18551\,
            in2 => \_gnd_net_\,
            in3 => \N__18560\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18536\,
            in2 => \_gnd_net_\,
            in3 => \N__18545\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19024\,
            in2 => \_gnd_net_\,
            in3 => \N__18530\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__19726\,
            in1 => \N__19169\,
            in2 => \_gnd_net_\,
            in3 => \N__18527\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19203\,
            in2 => \_gnd_net_\,
            in3 => \N__18524\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19252\,
            in2 => \_gnd_net_\,
            in3 => \N__18521\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19269\,
            in2 => \_gnd_net_\,
            in3 => \N__18518\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18981\,
            in2 => \_gnd_net_\,
            in3 => \N__18515\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19231\,
            in2 => \_gnd_net_\,
            in3 => \N__18611\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19182\,
            in2 => \_gnd_net_\,
            in3 => \N__18608\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19045\,
            in2 => \_gnd_net_\,
            in3 => \N__18605\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18602\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19300\,
            in2 => \_gnd_net_\,
            in3 => \N__19046\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19183\,
            in2 => \_gnd_net_\,
            in3 => \N__19327\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19369\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18983\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19396\,
            in2 => \_gnd_net_\,
            in3 => \N__19271\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18599\,
            in2 => \N__18587\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18839\,
            in2 => \N__18827\,
            in3 => \N__18815\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18812\,
            in2 => \N__18800\,
            in3 => \N__18788\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18785\,
            in2 => \N__18773\,
            in3 => \N__18761\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18758\,
            in2 => \N__18746\,
            in3 => \N__18728\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18725\,
            in2 => \N__18713\,
            in3 => \N__18698\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18695\,
            in2 => \N__18683\,
            in3 => \N__18668\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18665\,
            in2 => \N__18653\,
            in3 => \N__18638\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18635\,
            in2 => \N__18623\,
            in3 => \N__18614\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18965\,
            in2 => \N__18953\,
            in3 => \N__18941\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18938\,
            in2 => \N__19124\,
            in3 => \N__18926\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19112\,
            in2 => \N__18923\,
            in3 => \N__18908\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18905\,
            in2 => \N__19125\,
            in3 => \N__18893\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19116\,
            in2 => \N__18890\,
            in3 => \N__18875\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18872\,
            in2 => \N__19126\,
            in3 => \N__18860\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19120\,
            in2 => \N__18857\,
            in3 => \N__18845\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19517\,
            in1 => \N__19064\,
            in2 => \_gnd_net_\,
            in3 => \N__18842\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__19145\,
            in1 => \N__19105\,
            in2 => \N__20069\,
            in3 => \N__19076\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__20667\,
            in1 => \N__21264\,
            in2 => \N__20813\,
            in3 => \N__20520\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46103\,
            ce => 'H',
            sr => \N__45641\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__21265\,
            in1 => \N__20759\,
            in2 => \N__20522\,
            in3 => \N__20668\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46103\,
            ce => 'H',
            sr => \N__45641\
        );

    \rgb_drv_RNO_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__45726\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40576\,
            lcout => \rgb_drv_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_0_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__45727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40580\,
            lcout => \N_38_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__19044\,
            in1 => \N__19304\,
            in2 => \N__19760\,
            in3 => \N__19031\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19025\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19012\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__19013\,
            in1 => \N__18998\,
            in2 => \N__18992\,
            in3 => \N__19748\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__19749\,
            in1 => \N__18989\,
            in2 => \N__19376\,
            in3 => \N__18982\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__19277\,
            in1 => \N__19270\,
            in2 => \N__19400\,
            in3 => \N__19719\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19253\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19423\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__19424\,
            in1 => \N__19241\,
            in2 => \N__19235\,
            in3 => \N__19718\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19205\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19447\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19345\,
            in2 => \_gnd_net_\,
            in3 => \N__19232\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__19346\,
            in1 => \N__19220\,
            in2 => \N__19214\,
            in3 => \N__19754\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__19211\,
            in1 => \N__19204\,
            in2 => \N__19451\,
            in3 => \N__19717\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__19190\,
            in1 => \N__19184\,
            in2 => \N__19744\,
            in3 => \N__19328\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19168\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19463\,
            in2 => \_gnd_net_\,
            in3 => \N__19439\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19436\,
            in2 => \_gnd_net_\,
            in3 => \N__19415\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19412\,
            in2 => \_gnd_net_\,
            in3 => \N__19385\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19382\,
            in2 => \_gnd_net_\,
            in3 => \N__19358\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37669\,
            in2 => \N__19355\,
            in3 => \N__19337\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19334\,
            in2 => \N__37722\,
            in3 => \N__19316\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37673\,
            in2 => \N__19313\,
            in3 => \N__19289\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19286\,
            in2 => \_gnd_net_\,
            in3 => \N__19280\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19511\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19505\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19499\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19493\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19487\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19481\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19475\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19469\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19538\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19532\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19526\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19520\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21032\,
            in2 => \_gnd_net_\,
            in3 => \N__21053\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_5_LC_3_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19640\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46117\,
            ce => 'H',
            sr => \N__45579\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__20123\,
            in1 => \N__20064\,
            in2 => \N__19592\,
            in3 => \N__20270\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46115\,
            ce => 'H',
            sr => \N__45584\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__20273\,
            in1 => \N__20126\,
            in2 => \N__20077\,
            in3 => \N__19805\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46115\,
            ce => 'H',
            sr => \N__45584\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__20121\,
            in1 => \N__20062\,
            in2 => \N__19628\,
            in3 => \N__20268\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46115\,
            ce => 'H',
            sr => \N__45584\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_3_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__20124\,
            in1 => \N__20065\,
            in2 => \N__19574\,
            in3 => \N__20271\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46115\,
            ce => 'H',
            sr => \N__45584\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__20272\,
            in1 => \N__20125\,
            in2 => \N__20076\,
            in3 => \N__19547\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46115\,
            ce => 'H',
            sr => \N__45584\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__20122\,
            in1 => \N__20063\,
            in2 => \N__19610\,
            in3 => \N__20269\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46115\,
            ce => 'H',
            sr => \N__45584\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19634\,
            in2 => \N__19759\,
            in3 => \N__19753\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_8_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19619\,
            in2 => \_gnd_net_\,
            in3 => \N__19601\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19598\,
            in2 => \_gnd_net_\,
            in3 => \N__19583\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19580\,
            in2 => \_gnd_net_\,
            in3 => \N__19565\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19562\,
            in2 => \_gnd_net_\,
            in3 => \N__19556\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19553\,
            in2 => \_gnd_net_\,
            in3 => \N__19541\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19811\,
            in2 => \_gnd_net_\,
            in3 => \N__19799\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19796\,
            in2 => \_gnd_net_\,
            in3 => \N__19790\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19787\,
            in2 => \_gnd_net_\,
            in3 => \N__19781\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__19778\,
            in1 => \N__19769\,
            in2 => \N__19758\,
            in3 => \N__19667\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19654\,
            in1 => \N__19882\,
            in2 => \_gnd_net_\,
            in3 => \N__19909\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_duty_inputlt3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111011"
        )
    port map (
            in0 => \N__19865\,
            in1 => \N__20349\,
            in2 => \N__19664\,
            in3 => \N__20329\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__21277\,
            in1 => \N__20848\,
            in2 => \_gnd_net_\,
            in3 => \N__20196\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110010"
        )
    port map (
            in0 => \N__19921\,
            in1 => \N__20869\,
            in2 => \N__19853\,
            in3 => \N__20661\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__19849\,
            in1 => \N__20579\,
            in2 => \N__19661\,
            in3 => \N__19821\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46109\,
            ce => 'H',
            sr => \N__45602\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111111001101"
        )
    port map (
            in0 => \N__19922\,
            in1 => \N__20870\,
            in2 => \N__19855\,
            in3 => \N__20662\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46109\,
            ce => 'H',
            sr => \N__45602\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__19894\,
            in1 => \N__20558\,
            in2 => \N__19856\,
            in3 => \N__19823\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46109\,
            ce => 'H',
            sr => \N__45602\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__19822\,
            in1 => \N__20570\,
            in2 => \N__19854\,
            in3 => \N__19895\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46109\,
            ce => 'H',
            sr => \N__45602\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20428\,
            in2 => \_gnd_net_\,
            in3 => \N__20296\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__20373\,
            in1 => \N__20451\,
            in2 => \N__19868\,
            in3 => \N__20397\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__21269\,
            in1 => \N__20227\,
            in2 => \N__20216\,
            in3 => \N__20495\,
            lcout => \current_shift_inst.PI_CTRL.N_153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__20669\,
            in1 => \N__21270\,
            in2 => \_gnd_net_\,
            in3 => \N__20206\,
            lcout => \current_shift_inst.PI_CTRL.N_154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__20183\,
            in1 => \N__20849\,
            in2 => \N__20231\,
            in3 => \N__20506\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46099\,
            ce => 'H',
            sr => \N__45624\
        );

    \pwm_generator_inst.threshold_7_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20147\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46116\,
            ce => 'H',
            sr => \N__45574\
        );

    \pwm_generator_inst.threshold_2_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20177\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46116\,
            ce => 'H',
            sr => \N__45574\
        );

    \pwm_generator_inst.threshold_8_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46113\,
            ce => 'H',
            sr => \N__45580\
        );

    \pwm_generator_inst.threshold_3_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20171\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46113\,
            ce => 'H',
            sr => \N__45580\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__20117\,
            in1 => \N__20074\,
            in2 => \N__20165\,
            in3 => \N__20264\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46112\,
            ce => 'H',
            sr => \N__45585\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__20118\,
            in1 => \N__20075\,
            in2 => \N__20156\,
            in3 => \N__20265\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46112\,
            ce => 'H',
            sr => \N__45585\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__20266\,
            in1 => \N__20119\,
            in2 => \N__20078\,
            in3 => \N__20138\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46112\,
            ce => 'H',
            sr => \N__45585\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__20120\,
            in1 => \N__20267\,
            in2 => \N__20087\,
            in3 => \N__20073\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46112\,
            ce => 'H',
            sr => \N__45585\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20704\,
            in2 => \_gnd_net_\,
            in3 => \N__20802\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__20731\,
            in1 => \N__20752\,
            in2 => \N__19925\,
            in3 => \N__20779\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__21271\,
            in1 => \N__20665\,
            in2 => \N__20783\,
            in3 => \N__20515\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46104\,
            ce => 'H',
            sr => \N__45596\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100100010"
        )
    port map (
            in0 => \N__20664\,
            in1 => \N__21273\,
            in2 => \N__20521\,
            in3 => \N__20705\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46104\,
            ce => 'H',
            sr => \N__45596\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__21272\,
            in1 => \N__20666\,
            in2 => \N__20732\,
            in3 => \N__20516\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46104\,
            ce => 'H',
            sr => \N__45596\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20452\,
            in1 => \N__20432\,
            in2 => \N__20404\,
            in3 => \N__20374\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__20350\,
            in1 => \N__20330\,
            in2 => \N__20303\,
            in3 => \N__20300\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20697\,
            in2 => \_gnd_net_\,
            in3 => \N__20778\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20803\,
            in1 => \N__20751\,
            in2 => \N__20234\,
            in3 => \N__20727\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20834\,
            in2 => \_gnd_net_\,
            in3 => \N__20863\,
            lcout => \current_shift_inst.PI_CTRL.N_155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__21253\,
            in1 => \N__20835\,
            in2 => \N__20207\,
            in3 => \N__20663\,
            lcout => \current_shift_inst.PI_CTRL.N_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21139\,
            in1 => \N__20615\,
            in2 => \N__21314\,
            in3 => \N__20546\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20987\,
            in1 => \N__20975\,
            in2 => \N__20888\,
            in3 => \N__21065\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21121\,
            in2 => \_gnd_net_\,
            in3 => \N__21169\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21202\,
            in2 => \_gnd_net_\,
            in3 => \N__21187\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20974\,
            in1 => \N__20986\,
            in2 => \N__20540\,
            in3 => \N__21025\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20938\,
            in1 => \N__20887\,
            in2 => \N__20921\,
            in3 => \N__21064\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20477\,
            in1 => \N__20537\,
            in2 => \N__20531\,
            in3 => \N__20528\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20962\,
            in1 => \N__21082\,
            in2 => \N__21104\,
            in3 => \N__21292\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21293\,
            in1 => \N__20963\,
            in2 => \N__20471\,
            in3 => \N__21313\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20678\,
            in1 => \N__20609\,
            in2 => \N__20672\,
            in3 => \N__21110\,
            lcout => \current_shift_inst.PI_CTRL.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20998\,
            in1 => \N__21010\,
            in2 => \N__21158\,
            in3 => \N__21046\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21011\,
            in1 => \N__20999\,
            in2 => \N__20945\,
            in3 => \N__20920\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23664\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21385\,
            ce => 'H',
            sr => \N__45654\
        );

    \pwm_generator_inst.threshold_1_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20603\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46114\,
            ce => 'H',
            sr => \N__45568\
        );

    \pwm_generator_inst.threshold_0_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20591\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46114\,
            ce => 'H',
            sr => \N__45568\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21416\,
            in2 => \N__24125\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__46100\,
            ce => 'H',
            sr => \N__45591\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21407\,
            in2 => \N__26414\,
            in3 => \N__20561\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__46100\,
            ce => 'H',
            sr => \N__45591\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21584\,
            in2 => \N__24053\,
            in3 => \N__20549\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__46100\,
            ce => 'H',
            sr => \N__45591\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21791\,
            in2 => \N__23981\,
            in3 => \N__20852\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__46100\,
            ce => 'H',
            sr => \N__45591\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21575\,
            in2 => \N__22907\,
            in3 => \N__20816\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__46100\,
            ce => 'H',
            sr => \N__45591\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21566\,
            in2 => \N__26153\,
            in3 => \N__20786\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__46100\,
            ce => 'H',
            sr => \N__45591\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21539\,
            in2 => \N__27530\,
            in3 => \N__20762\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__46100\,
            ce => 'H',
            sr => \N__45591\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21593\,
            in2 => \N__22319\,
            in3 => \N__20735\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__46100\,
            ce => 'H',
            sr => \N__45591\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23882\,
            in2 => \N__21398\,
            in3 => \N__20708\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__46095\,
            ce => 'H',
            sr => \N__45597\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21425\,
            in2 => \N__24194\,
            in3 => \N__20684\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__46095\,
            ce => 'H',
            sr => \N__45597\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21548\,
            in2 => \N__26942\,
            in3 => \N__20681\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__46095\,
            ce => 'H',
            sr => \N__45597\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21557\,
            in2 => \N__22661\,
            in3 => \N__20951\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__46095\,
            ce => 'H',
            sr => \N__45597\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21447\,
            in2 => \N__22505\,
            in3 => \N__20948\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__46095\,
            ce => 'H',
            sr => \N__45597\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22742\,
            in2 => \N__21489\,
            in3 => \N__20924\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__46095\,
            ce => 'H',
            sr => \N__45597\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21451\,
            in2 => \N__26342\,
            in3 => \N__20903\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__46095\,
            ce => 'H',
            sr => \N__45597\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23144\,
            in2 => \N__21490\,
            in3 => \N__20900\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__46095\,
            ce => 'H',
            sr => \N__45597\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21491\,
            in2 => \N__23294\,
            in3 => \N__20897\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__46089\,
            ce => 'H',
            sr => \N__45603\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23234\,
            in2 => \N__21521\,
            in3 => \N__20894\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__46089\,
            ce => 'H',
            sr => \N__45603\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21495\,
            in2 => \N__22994\,
            in3 => \N__20891\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__46089\,
            ce => 'H',
            sr => \N__45603\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26288\,
            in2 => \N__21522\,
            in3 => \N__20873\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__46089\,
            ce => 'H',
            sr => \N__45603\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21499\,
            in2 => \N__26819\,
            in3 => \N__21056\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__46089\,
            ce => 'H',
            sr => \N__45603\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26563\,
            in2 => \N__21523\,
            in3 => \N__21035\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__46089\,
            ce => 'H',
            sr => \N__45603\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21503\,
            in2 => \N__26687\,
            in3 => \N__21014\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__46089\,
            ce => 'H',
            sr => \N__45603\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24882\,
            in2 => \N__21524\,
            in3 => \N__21002\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__46089\,
            ce => 'H',
            sr => \N__45603\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21507\,
            in2 => \N__23522\,
            in3 => \N__20990\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__46080\,
            ce => 'H',
            sr => \N__45611\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23428\,
            in2 => \N__21525\,
            in3 => \N__20978\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__46080\,
            ce => 'H',
            sr => \N__45611\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21511\,
            in2 => \N__23374\,
            in3 => \N__20966\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__46080\,
            ce => 'H',
            sr => \N__45611\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31408\,
            in2 => \N__21526\,
            in3 => \N__20954\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__46080\,
            ce => 'H',
            sr => \N__45611\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21515\,
            in2 => \N__31352\,
            in3 => \N__21299\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__46080\,
            ce => 'H',
            sr => \N__45611\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27464\,
            in2 => \N__21527\,
            in3 => \N__21296\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__46080\,
            ce => 'H',
            sr => \N__45611\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21519\,
            in2 => \N__31463\,
            in3 => \N__21284\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__46080\,
            ce => 'H',
            sr => \N__45611\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21520\,
            in1 => \N__27404\,
            in2 => \_gnd_net_\,
            in3 => \N__21281\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46080\,
            ce => 'H',
            sr => \N__45611\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21206\,
            in1 => \N__21191\,
            in2 => \N__21176\,
            in3 => \N__21157\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21143\,
            in1 => \N__21071\,
            in2 => \N__21128\,
            in3 => \N__21125\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24049\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21100\,
            in2 => \_gnd_net_\,
            in3 => \N__21086\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36917\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46068\,
            ce => 'H',
            sr => \N__45633\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21913\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46068\,
            ce => 'H',
            sr => \N__45633\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21893\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46068\,
            ce => 'H',
            sr => \N__45633\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22861\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46068\,
            ce => 'H',
            sr => \N__45633\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31610\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46042\,
            ce => \N__33768\,
            sr => \N__45652\
        );

    \delay_measurement_inst.stop_timer_hc_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23665\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21386\,
            ce => 'H',
            sr => \N__45655\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21374\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_6_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21347\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46110\,
            ce => 'H',
            sr => \N__45561\
        );

    \pwm_generator_inst.threshold_4_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21335\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46105\,
            ce => 'H',
            sr => \N__45565\
        );

    \pwm_generator_inst.threshold_9_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21323\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46101\,
            ce => 'H',
            sr => \N__45569\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26462\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46090\,
            ce => 'H',
            sr => \N__45581\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21872\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46090\,
            ce => 'H',
            sr => \N__45581\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26758\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46090\,
            ce => 'H',
            sr => \N__45581\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22816\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46090\,
            ce => 'H',
            sr => \N__45581\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21815\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46081\,
            ce => 'H',
            sr => \N__45586\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27587\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46081\,
            ce => 'H',
            sr => \N__45586\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22444\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46081\,
            ce => 'H',
            sr => \N__45586\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33047\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46081\,
            ce => 'H',
            sr => \N__45586\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26212\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46081\,
            ce => 'H',
            sr => \N__45586\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23417\,
            in1 => \N__31391\,
            in2 => \N__31345\,
            in3 => \N__23361\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21605\,
            in1 => \N__22589\,
            in2 => \N__21608\,
            in3 => \N__21758\,
            lcout => \current_shift_inst.PI_CTRL.N_74_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26679\,
            in1 => \N__23511\,
            in2 => \N__26564\,
            in3 => \N__26283\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31338\,
            in2 => \_gnd_net_\,
            in3 => \N__23416\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31459\,
            in1 => \N__31390\,
            in2 => \N__21599\,
            in3 => \N__21614\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__26149\,
            in1 => \N__22906\,
            in2 => \N__23980\,
            in3 => \N__22277\,
            lcout => \current_shift_inst.PI_CTRL.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23138\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22975\,
            in1 => \N__23223\,
            in2 => \N__23139\,
            in3 => \N__26811\,
            lcout => \current_shift_inst.PI_CTRL.N_74_16\,
            ltout => \current_shift_inst.PI_CTRL.N_74_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21625\,
            in1 => \N__21634\,
            in2 => \N__21596\,
            in3 => \N__22649\,
            lcout => \current_shift_inst.PI_CTRL.N_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26138\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36899\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23501\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27395\,
            in1 => \N__21641\,
            in2 => \_gnd_net_\,
            in3 => \N__22648\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__21635\,
            in1 => \N__21626\,
            in2 => \N__21617\,
            in3 => \N__21770\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23500\,
            in1 => \N__26273\,
            in2 => \N__26559\,
            in3 => \N__23347\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__27193\,
            in1 => \N__27398\,
            in2 => \N__24209\,
            in3 => \N__27035\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46062\,
            ce => 'H',
            sr => \N__45604\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22638\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__27396\,
            in1 => \N__27196\,
            in2 => \N__27090\,
            in3 => \N__24776\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46062\,
            ce => 'H',
            sr => \N__45604\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__27194\,
            in1 => \N__27399\,
            in2 => \N__24737\,
            in3 => \N__27036\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46062\,
            ce => 'H',
            sr => \N__45604\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__27397\,
            in1 => \N__27197\,
            in2 => \N__27091\,
            in3 => \N__24698\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46062\,
            ce => 'H',
            sr => \N__45604\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__27195\,
            in1 => \N__27400\,
            in2 => \N__24659\,
            in3 => \N__27037\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46062\,
            ce => 'H',
            sr => \N__45604\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21674\,
            in2 => \_gnd_net_\,
            in3 => \N__36916\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21668\,
            in2 => \_gnd_net_\,
            in3 => \N__21659\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45612\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26228\,
            in2 => \_gnd_net_\,
            in3 => \N__21656\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45612\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26720\,
            in2 => \_gnd_net_\,
            in3 => \N__21653\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45612\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22073\,
            in2 => \_gnd_net_\,
            in3 => \N__21650\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45612\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23162\,
            in2 => \_gnd_net_\,
            in3 => \N__21647\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45612\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26828\,
            in2 => \_gnd_net_\,
            in3 => \N__21644\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45612\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21824\,
            in2 => \_gnd_net_\,
            in3 => \N__21692\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45612\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33158\,
            in2 => \_gnd_net_\,
            in3 => \N__21689\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__46048\,
            ce => 'H',
            sr => \N__45625\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47387\,
            in2 => \_gnd_net_\,
            in3 => \N__21686\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__46048\,
            ce => 'H',
            sr => \N__45625\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31628\,
            in2 => \_gnd_net_\,
            in3 => \N__21683\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__46048\,
            ce => 'H',
            sr => \N__45625\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36998\,
            in2 => \_gnd_net_\,
            in3 => \N__21680\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__46048\,
            ce => 'H',
            sr => \N__45625\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37037\,
            in2 => \_gnd_net_\,
            in3 => \N__21677\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46048\,
            ce => 'H',
            sr => \N__45625\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22845\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26202\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27579\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22525\,
            in2 => \_gnd_net_\,
            in3 => \N__32943\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22939\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23092\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32946\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32944\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22705\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23479\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32950\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32945\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22558\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__24826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32949\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32947\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23314\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__23813\,
            in1 => \N__23599\,
            in2 => \N__28494\,
            in3 => \N__22046\,
            lcout => \phase_controller_inst1.stoper_hc.N_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__28242\,
            in1 => \N__23576\,
            in2 => \N__27878\,
            in3 => \N__23600\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46036\,
            ce => \N__28873\,
            sr => \N__45637\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101110"
        )
    port map (
            in0 => \N__23605\,
            in1 => \N__30202\,
            in2 => \N__30485\,
            in3 => \N__41565\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__23769\,
            in1 => \N__41567\,
            in2 => \N__30701\,
            in3 => \N__30204\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21746\,
            in3 => \N__30270\,
            lcout => \elapsed_time_ns_1_RNI51CED1_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__23827\,
            in1 => \N__41566\,
            in2 => \N__30347\,
            in3 => \N__30203\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23031\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33046\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100100"
        )
    port map (
            in0 => \N__41569\,
            in1 => \N__23712\,
            in2 => \N__30665\,
            in3 => \N__30206\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28685\,
            in2 => \_gnd_net_\,
            in3 => \N__23640\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_432_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21728\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21719\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21704\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46091\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21851\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46082\,
            ce => 'H',
            sr => \N__45575\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21814\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__22650\,
            in1 => \N__26680\,
            in2 => \_gnd_net_\,
            in3 => \N__21752\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22397\,
            in1 => \N__22403\,
            in2 => \N__21782\,
            in3 => \N__21779\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__21764\,
            in1 => \N__22895\,
            in2 => \N__21773\,
            in3 => \N__22409\,
            lcout => \current_shift_inst.PI_CTRL.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111111111"
        )
    port map (
            in0 => \N__24048\,
            in1 => \N__26410\,
            in2 => \N__24124\,
            in3 => \N__23973\,
            lcout => \current_shift_inst.PI_CTRL.N_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23360\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24881\,
            in1 => \N__27459\,
            in2 => \N__23289\,
            in3 => \N__26937\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__22770\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33048\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26803\,
            in1 => \N__23221\,
            in2 => \N__22985\,
            in3 => \N__23128\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22440\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37097\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26637\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23266\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23959\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24111\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__22298\,
            in1 => \N__21813\,
            in2 => \N__33131\,
            in3 => \N__21932\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22297\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__27200\,
            in1 => \N__27391\,
            in2 => \N__27094\,
            in3 => \N__24320\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46055\,
            ce => 'H',
            sr => \N__45598\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__27387\,
            in1 => \N__27201\,
            in2 => \N__24515\,
            in3 => \N__27047\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46055\,
            ce => 'H',
            sr => \N__45598\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__27198\,
            in1 => \N__27389\,
            in2 => \N__27092\,
            in3 => \N__24470\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46055\,
            ce => 'H',
            sr => \N__45598\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__27388\,
            in1 => \N__27202\,
            in2 => \N__24440\,
            in3 => \N__27048\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46055\,
            ce => 'H',
            sr => \N__45598\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__27199\,
            in1 => \N__27390\,
            in2 => \N__27093\,
            in3 => \N__24398\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46055\,
            ce => 'H',
            sr => \N__45598\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21899\,
            in2 => \_gnd_net_\,
            in3 => \N__21914\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21878\,
            in2 => \_gnd_net_\,
            in3 => \N__21889\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21857\,
            in2 => \_gnd_net_\,
            in3 => \N__21868\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21833\,
            in2 => \_gnd_net_\,
            in3 => \N__21844\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26729\,
            in2 => \_gnd_net_\,
            in3 => \N__21827\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22787\,
            in2 => \_gnd_net_\,
            in3 => \N__21986\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21983\,
            in2 => \_gnd_net_\,
            in3 => \N__21974\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26426\,
            in2 => \_gnd_net_\,
            in3 => \N__21971\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21968\,
            in2 => \_gnd_net_\,
            in3 => \N__21962\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_8\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21959\,
            in2 => \_gnd_net_\,
            in3 => \N__21953\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21950\,
            in2 => \_gnd_net_\,
            in3 => \N__21944\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21941\,
            in2 => \_gnd_net_\,
            in3 => \N__21923\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23061\,
            in2 => \_gnd_net_\,
            in3 => \N__21920\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23010\,
            in2 => \_gnd_net_\,
            in3 => \N__21917\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22771\,
            in2 => \_gnd_net_\,
            in3 => \N__22013\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22672\,
            in2 => \_gnd_net_\,
            in3 => \N__22010\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22521\,
            in2 => \_gnd_net_\,
            in3 => \N__22007\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22695\,
            in2 => \_gnd_net_\,
            in3 => \N__22004\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22554\,
            in2 => \_gnd_net_\,
            in3 => \N__22001\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23088\,
            in2 => \_gnd_net_\,
            in3 => \N__21998\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23310\,
            in2 => \_gnd_net_\,
            in3 => \N__21995\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23194\,
            in2 => \_gnd_net_\,
            in3 => \N__21992\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22935\,
            in2 => \_gnd_net_\,
            in3 => \N__21989\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26710\,
            in2 => \_gnd_net_\,
            in3 => \N__22040\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23032\,
            in2 => \_gnd_net_\,
            in3 => \N__22037\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26593\,
            in2 => \_gnd_net_\,
            in3 => \N__22034\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26638\,
            in2 => \_gnd_net_\,
            in3 => \N__22031\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24822\,
            in2 => \_gnd_net_\,
            in3 => \N__22028\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23475\,
            in2 => \_gnd_net_\,
            in3 => \N__22025\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23452\,
            in2 => \_gnd_net_\,
            in3 => \N__22022\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23386\,
            in2 => \_gnd_net_\,
            in3 => \N__22019\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__33111\,
            in1 => \N__31409\,
            in2 => \_gnd_net_\,
            in3 => \N__22016\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22079\,
            in2 => \_gnd_net_\,
            in3 => \N__30265\,
            lcout => \elapsed_time_ns_1_RNIL13KD1_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37148\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__22061\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30266\,
            lcout => \elapsed_time_ns_1_RNI1TBED1_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111101100"
        )
    port map (
            in0 => \N__41545\,
            in1 => \N__30200\,
            in2 => \N__30767\,
            in3 => \N__23549\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22055\,
            in3 => \N__30264\,
            lcout => \elapsed_time_ns_1_RNI3VBED1_0_16\,
            ltout => \elapsed_time_ns_1_RNI3VBED1_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28339\,
            in1 => \N__23732\,
            in2 => \N__22052\,
            in3 => \N__28086\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23708\,
            in2 => \N__22049\,
            in3 => \N__23762\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__23763\,
            in1 => \N__23550\,
            in2 => \N__23714\,
            in3 => \N__23742\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22130\,
            in2 => \_gnd_net_\,
            in3 => \N__30263\,
            lcout => \elapsed_time_ns_1_RNI40CED1_0_17\,
            ltout => \elapsed_time_ns_1_RNI40CED1_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010111010"
        )
    port map (
            in0 => \N__30205\,
            in1 => \N__41568\,
            in2 => \N__22133\,
            in3 => \N__30731\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_14_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28481\,
            in2 => \_gnd_net_\,
            in3 => \N__27752\,
            lcout => \phase_controller_inst1.stoper_hc.N_287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__45723\,
            in1 => \N__27992\,
            in2 => \N__28564\,
            in3 => \N__29900\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__28603\,
            in1 => \_gnd_net_\,
            in2 => \N__22124\,
            in3 => \N__29930\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__45722\,
            in1 => \N__28604\,
            in2 => \N__28565\,
            in3 => \N__29876\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__45724\,
            in1 => \N__30850\,
            in2 => \N__22121\,
            in3 => \N__22118\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__22112\,
            in1 => \_gnd_net_\,
            in2 => \N__22103\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNI62CED1_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__28489\,
            in1 => \N__23828\,
            in2 => \_gnd_net_\,
            in3 => \N__27751\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_8_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__28690\,
            in1 => \N__23678\,
            in2 => \_gnd_net_\,
            in3 => \N__23644\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46008\,
            ce => 'H',
            sr => \N__45657\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22100\,
            in2 => \N__22091\,
            in3 => \N__25682\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22268\,
            in2 => \N__22259\,
            in3 => \N__26075\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22250\,
            in2 => \N__22241\,
            in3 => \N__26048\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22232\,
            in2 => \N__22217\,
            in3 => \N__26024\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25997\,
            in1 => \N__22208\,
            in2 => \N__22196\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25973\,
            in1 => \N__22187\,
            in2 => \N__22178\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22157\,
            in2 => \N__22169\,
            in3 => \N__25949\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22139\,
            in2 => \N__22151\,
            in3 => \N__25922\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22391\,
            in2 => \N__22382\,
            in3 => \N__25898\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22373\,
            in2 => \N__22361\,
            in3 => \N__25832\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22352\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46096\,
            ce => 'H',
            sr => \N__45557\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22328\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22308\,
            in2 => \_gnd_net_\,
            in3 => \N__26142\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23427\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22990\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22318\,
            in1 => \N__23867\,
            in2 => \N__27528\,
            in3 => \N__24179\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22731\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__22415\,
            in1 => \N__23868\,
            in2 => \N__27529\,
            in3 => \N__24180\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24880\,
            in1 => \N__23279\,
            in2 => \N__26938\,
            in3 => \N__27458\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22486\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26586\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33049\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22888\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__27378\,
            in1 => \N__27224\,
            in2 => \N__27114\,
            in3 => \N__24371\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46056\,
            ce => 'H',
            sr => \N__45587\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__27221\,
            in1 => \N__27379\,
            in2 => \N__27115\,
            in3 => \N__24593\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46056\,
            ce => 'H',
            sr => \N__45587\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__27376\,
            in1 => \N__27222\,
            in2 => \N__27112\,
            in3 => \N__24566\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46056\,
            ce => 'H',
            sr => \N__45587\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26327\,
            in1 => \N__22729\,
            in2 => \N__22498\,
            in3 => \N__27375\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__27377\,
            in1 => \N__27223\,
            in2 => \N__27113\,
            in3 => \N__24548\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46056\,
            ce => 'H',
            sr => \N__45587\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26326\,
            in1 => \N__22730\,
            in2 => \N__22497\,
            in3 => \N__31455\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101111"
        )
    port map (
            in0 => \N__22577\,
            in1 => \N__24148\,
            in2 => \N__33128\,
            in3 => \N__26759\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__22571\,
            in1 => \N__26400\,
            in2 => \N__22820\,
            in3 => \N__33088\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__22565\,
            in1 => \N__26331\,
            in2 => \N__33130\,
            in3 => \N__22538\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23222\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__22529\,
            in1 => \N__22496\,
            in2 => \N__33129\,
            in3 => \N__22463\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__24038\,
            in1 => \N__22454\,
            in2 => \N__22448\,
            in3 => \N__33089\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27460\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__22896\,
            in1 => \N__33090\,
            in2 => \N__22862\,
            in3 => \N__22829\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22812\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__24190\,
            in1 => \N__23011\,
            in2 => \N__33126\,
            in3 => \N__22781\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__26930\,
            in1 => \N__33076\,
            in2 => \N__22775\,
            in3 => \N__22748\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__22741\,
            in1 => \N__22706\,
            in2 => \N__33127\,
            in3 => \N__22682\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22673\,
            in2 => \_gnd_net_\,
            in3 => \N__33073\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__33080\,
            in1 => \N__22660\,
            in2 => \N__22616\,
            in3 => \N__22613\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__26461\,
            in1 => \N__23969\,
            in2 => \N__22607\,
            in3 => \N__33074\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__33075\,
            in1 => \N__23878\,
            in2 => \N__23066\,
            in3 => \N__22595\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__23233\,
            in1 => \N__23195\,
            in2 => \N__33066\,
            in3 => \N__23171\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37127\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__26287\,
            in1 => \N__26711\,
            in2 => \N__33067\,
            in3 => \N__23150\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__23143\,
            in1 => \N__32978\,
            in2 => \N__23099\,
            in3 => \N__23072\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23065\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111101101111"
        )
    port map (
            in0 => \N__23045\,
            in1 => \N__23036\,
            in2 => \N__33132\,
            in3 => \N__26815\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__23012\,
            in1 => \_gnd_net_\,
            in2 => \N__33065\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011111111"
        )
    port map (
            in0 => \N__22989\,
            in1 => \N__22943\,
            in2 => \N__22919\,
            in3 => \N__32982\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__23521\,
            in1 => \N__23480\,
            in2 => \N__33133\,
            in3 => \N__23459\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23453\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33103\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110101111101"
        )
    port map (
            in0 => \N__33110\,
            in1 => \N__23441\,
            in2 => \N__23432\,
            in3 => \N__23429\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23387\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33104\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__33109\,
            in1 => \N__23375\,
            in2 => \N__23324\,
            in3 => \N__23321\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.N_266_i_1_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010000"
        )
    port map (
            in0 => \N__27753\,
            in1 => \N__24977\,
            in2 => \N__28496\,
            in3 => \N__23829\,
            lcout => \phase_controller_inst1.stoper_hc.N_266_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__23315\,
            in1 => \N__23290\,
            in2 => \N__23246\,
            in3 => \N__33105\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__23814\,
            in1 => \N__23601\,
            in2 => \_gnd_net_\,
            in3 => \N__24975\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.N_275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010000"
        )
    port map (
            in0 => \N__28485\,
            in1 => \N__27810\,
            in2 => \N__23237\,
            in3 => \N__27744\,
            lcout => \phase_controller_inst1.stoper_hc.N_325\,
            ltout => \phase_controller_inst1.stoper_hc.N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28173\,
            in2 => \N__23531\,
            in3 => \N__27628\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__27629\,
            in1 => \N__28064\,
            in2 => \N__23528\,
            in3 => \N__27599\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46031\,
            ce => \N__28872\,
            sr => \N__45626\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__28063\,
            in1 => \N__28175\,
            in2 => \N__28310\,
            in3 => \N__30233\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46031\,
            ce => \N__28872\,
            sr => \N__45626\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__28174\,
            in1 => \N__28065\,
            in2 => \N__28361\,
            in3 => \N__28298\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46031\,
            ce => \N__28872\,
            sr => \N__45626\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__28290\,
            in1 => \N__28068\,
            in2 => \N__28343\,
            in3 => \N__28228\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46027\,
            ce => \N__28871\,
            sr => \N__45634\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__41711\,
            in1 => \N__41544\,
            in2 => \N__30083\,
            in3 => \N__28090\,
            lcout => \elapsed_time_ns_1_RNIB4DJ11_0_5\,
            ltout => \elapsed_time_ns_1_RNIB4DJ11_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__28291\,
            in1 => \N__28069\,
            in2 => \N__23525\,
            in3 => \N__28229\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46027\,
            ce => \N__28871\,
            sr => \N__45634\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__28292\,
            in1 => \N__28227\,
            in2 => \_gnd_net_\,
            in3 => \N__27707\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46027\,
            ce => \N__28871\,
            sr => \N__45634\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__28226\,
            in1 => \N__27680\,
            in2 => \_gnd_net_\,
            in3 => \N__28294\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46027\,
            ce => \N__28871\,
            sr => \N__45634\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__28067\,
            in1 => \N__28649\,
            in2 => \N__27650\,
            in3 => \N__28293\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46027\,
            ce => \N__28871\,
            sr => \N__45634\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010001"
        )
    port map (
            in0 => \N__28233\,
            in1 => \N__23845\,
            in2 => \N__23833\,
            in3 => \N__27855\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46023\,
            ce => \N__29308\,
            sr => \N__45638\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__23707\,
            in1 => \N__27856\,
            in2 => \_gnd_net_\,
            in3 => \N__28236\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46023\,
            ce => \N__29308\,
            sr => \N__45638\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__28231\,
            in1 => \N__23776\,
            in2 => \_gnd_net_\,
            in3 => \N__27853\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46023\,
            ce => \N__29308\,
            sr => \N__45638\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__27850\,
            in1 => \N__28234\,
            in2 => \_gnd_net_\,
            in3 => \N__23744\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46023\,
            ce => \N__29308\,
            sr => \N__45638\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__28230\,
            in1 => \N__27852\,
            in2 => \_gnd_net_\,
            in3 => \N__23554\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46023\,
            ce => \N__29308\,
            sr => \N__45638\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__27851\,
            in1 => \N__28235\,
            in2 => \N__23606\,
            in3 => \N__23572\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46023\,
            ce => \N__29308\,
            sr => \N__45638\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__28232\,
            in1 => \N__25038\,
            in2 => \N__27957\,
            in3 => \N__27854\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46023\,
            ce => \N__29308\,
            sr => \N__45638\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__28243\,
            in1 => \N__27939\,
            in2 => \N__25046\,
            in3 => \N__27864\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46020\,
            ce => \N__28874\,
            sr => \N__45642\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__27861\,
            in1 => \N__28246\,
            in2 => \_gnd_net_\,
            in3 => \N__23555\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46020\,
            ce => \N__28874\,
            sr => \N__45642\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__27862\,
            in1 => \N__28247\,
            in2 => \N__27761\,
            in3 => \N__28490\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46020\,
            ce => \N__28874\,
            sr => \N__45642\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010001"
        )
    port map (
            in0 => \N__28245\,
            in1 => \N__23846\,
            in2 => \N__23834\,
            in3 => \N__27865\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46020\,
            ce => \N__28874\,
            sr => \N__45642\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__28244\,
            in1 => \N__27863\,
            in2 => \N__27964\,
            in3 => \N__26890\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46020\,
            ce => \N__28874\,
            sr => \N__45642\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27868\,
            in1 => \N__28241\,
            in2 => \N__26864\,
            in3 => \N__27946\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => \N__28862\,
            sr => \N__45649\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__28238\,
            in1 => \N__27908\,
            in2 => \N__27958\,
            in3 => \N__27870\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => \N__28862\,
            sr => \N__45649\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__27866\,
            in1 => \N__28239\,
            in2 => \_gnd_net_\,
            in3 => \N__23777\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => \N__28862\,
            sr => \N__45649\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__28237\,
            in1 => \N__27869\,
            in2 => \_gnd_net_\,
            in3 => \N__23743\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => \N__28862\,
            sr => \N__45649\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__27867\,
            in1 => \N__28240\,
            in2 => \_gnd_net_\,
            in3 => \N__23713\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => \N__28862\,
            sr => \N__45649\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__28689\,
            in1 => \N__23677\,
            in2 => \_gnd_net_\,
            in3 => \N__23645\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_433_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S1_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41982\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45992\,
            ce => 'H',
            sr => \N__45662\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25827\,
            in1 => \N__25893\,
            in2 => \_gnd_net_\,
            in3 => \N__25920\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26043\,
            in2 => \_gnd_net_\,
            in3 => \N__25677\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__25995\,
            in1 => \N__26019\,
            in2 => \N__23912\,
            in3 => \N__26073\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23909\,
            in1 => \N__25944\,
            in2 => \N__23903\,
            in3 => \N__25972\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23900\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23888\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31074\,
            in2 => \_gnd_net_\,
            in3 => \N__29097\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23866\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__27238\,
            in1 => \N__27403\,
            in2 => \N__27116\,
            in3 => \N__24290\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46050\,
            ce => 'H',
            sr => \N__45570\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__27402\,
            in1 => \N__27240\,
            in2 => \N__24257\,
            in3 => \N__27099\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46050\,
            ce => 'H',
            sr => \N__45570\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24167\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__27401\,
            in1 => \N__27239\,
            in2 => \N__24626\,
            in3 => \N__27098\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46050\,
            ce => 'H',
            sr => \N__45570\
        );

    \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26353\,
            in2 => \N__26357\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__27088\,
            in1 => \N__24149\,
            in2 => \N__24134\,
            in3 => \N__24089\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            clk => \N__46044\,
            ce => 'H',
            sr => \N__45576\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__27069\,
            in1 => \N__24086\,
            in2 => \N__26372\,
            in3 => \N__24080\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            clk => \N__46044\,
            ce => 'H',
            sr => \N__45576\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__27089\,
            in1 => \N__24077\,
            in2 => \N__24062\,
            in3 => \N__24005\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            clk => \N__46044\,
            ce => 'H',
            sr => \N__45576\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0111110111010111"
        )
    port map (
            in0 => \N__27070\,
            in1 => \N__24002\,
            in2 => \N__23993\,
            in3 => \N__23930\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            clk => \N__46044\,
            ce => 'H',
            sr => \N__45576\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23927\,
            in2 => \N__23921\,
            in3 => \N__24365\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24362\,
            in2 => \N__26174\,
            in3 => \N__24350\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26237\,
            in2 => \N__27554\,
            in3 => \N__24347\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24344\,
            in2 => \N__24335\,
            in3 => \N__24311\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24308\,
            in2 => \N__24299\,
            in3 => \N__24281\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24278\,
            in2 => \N__24266\,
            in3 => \N__24245\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26834\,
            in2 => \N__24242\,
            in3 => \N__24230\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24227\,
            in2 => \N__24218\,
            in3 => \N__24197\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24611\,
            in2 => \N__24602\,
            in3 => \N__24587\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24584\,
            in2 => \N__24575\,
            in3 => \N__24560\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26300\,
            in2 => \N__24557\,
            in3 => \N__24542\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24539\,
            in2 => \N__24527\,
            in3 => \N__24500\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24497\,
            in2 => \N__24485\,
            in3 => \N__24458\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24455\,
            in2 => \N__24449\,
            in3 => \N__24422\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24419\,
            in2 => \N__24407\,
            in3 => \N__24386\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26243\,
            in2 => \N__24383\,
            in3 => \N__24374\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26768\,
            in2 => \N__24794\,
            in3 => \N__24785\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26363\,
            in2 => \N__26495\,
            in3 => \N__24782\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26294\,
            in2 => \N__26603\,
            in3 => \N__24779\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24890\,
            in2 => \N__24806\,
            in3 => \N__24764\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24761\,
            in2 => \N__24749\,
            in3 => \N__24722\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24719\,
            in2 => \N__24707\,
            in3 => \N__24686\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24683\,
            in2 => \N__24671\,
            in3 => \N__24644\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31361\,
            in2 => \N__24641\,
            in3 => \N__24614\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31307\,
            in2 => \N__32857\,
            in3 => \N__24914\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32853\,
            in2 => \N__24911\,
            in3 => \N__24899\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31418\,
            in2 => \N__32858\,
            in3 => \N__24896\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__33136\,
            in1 => \N__27310\,
            in2 => \_gnd_net_\,
            in3 => \N__24893\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__41716\,
            in1 => \N__41575\,
            in2 => \N__30512\,
            in3 => \N__27678\,
            lcout => \elapsed_time_ns_1_RNIE7DJ11_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24883\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__47048\,
            in1 => \N__47337\,
            in2 => \N__46397\,
            in3 => \N__47002\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__33135\,
            in1 => \N__24884\,
            in2 => \N__24842\,
            in3 => \N__24827\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110011"
        )
    port map (
            in0 => \N__28644\,
            in1 => \N__41387\,
            in2 => \N__24944\,
            in3 => \N__24959\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__41715\,
            in1 => \N__41574\,
            in2 => \N__30539\,
            in3 => \N__27706\,
            lcout => \elapsed_time_ns_1_RNID6DJ11_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__27701\,
            in1 => \N__24976\,
            in2 => \N__27679\,
            in3 => \N__30232\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__28480\,
            in1 => \_gnd_net_\,
            in2 => \N__24983\,
            in3 => \N__27811\,
            lcout => \phase_controller_inst1.stoper_hc.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__41519\,
            in1 => \N__41702\,
            in2 => \N__30371\,
            in3 => \N__27897\,
            lcout => \elapsed_time_ns_1_RNIQ2MD11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__26847\,
            in1 => \N__41518\,
            in2 => \N__30395\,
            in3 => \N__41700\,
            lcout => \elapsed_time_ns_1_RNIP1MD11_0_12\,
            ltout => \elapsed_time_ns_1_RNIP1MD11_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25031\,
            in1 => \N__27896\,
            in2 => \N__24980\,
            in3 => \N__26882\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__24958\,
            in1 => \N__28176\,
            in2 => \N__24943\,
            in3 => \N__27815\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__28613\,
            in1 => \N__24957\,
            in2 => \N__27857\,
            in3 => \N__24939\,
            lcout => \phase_controller_inst1.stoper_hc.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__26883\,
            in1 => \N__41701\,
            in2 => \N__30419\,
            in3 => \N__41520\,
            lcout => \elapsed_time_ns_1_RNIO0MD11_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__41497\,
            in1 => \N__41692\,
            in2 => \N__30446\,
            in3 => \N__25042\,
            lcout => \elapsed_time_ns_1_RNINVLD11_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__41689\,
            in1 => \N__41496\,
            in2 => \N__30107\,
            in3 => \N__28338\,
            lcout => \elapsed_time_ns_1_RNIA3DJ11_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__41498\,
            in1 => \N__25013\,
            in2 => \N__30608\,
            in3 => \N__41691\,
            lcout => \elapsed_time_ns_1_RNIP2ND11_0_21\,
            ltout => \elapsed_time_ns_1_RNIP2ND11_0_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25000\,
            in1 => \N__28507\,
            in2 => \N__25007\,
            in3 => \N__28393\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25124\,
            in1 => \N__25142\,
            in2 => \N__25004\,
            in3 => \N__25108\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__28007\,
            in1 => \N__29929\,
            in2 => \N__27991\,
            in3 => \N__30854\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__41499\,
            in1 => \N__41693\,
            in2 => \N__30971\,
            in3 => \N__25001\,
            lcout => \elapsed_time_ns_1_RNIU7ND11_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41690\,
            in1 => \N__25136\,
            in2 => \N__41550\,
            in3 => \N__30926\,
            lcout => \elapsed_time_ns_1_RNI0AND11_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__24992\,
            in1 => \N__41688\,
            in2 => \N__30566\,
            in3 => \N__41500\,
            lcout => \elapsed_time_ns_1_RNIR4ND11_0_23\,
            ltout => \elapsed_time_ns_1_RNIR4ND11_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28018\,
            in1 => \N__28519\,
            in2 => \N__24986\,
            in3 => \N__25117\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25135\,
            in2 => \_gnd_net_\,
            in3 => \N__25093\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__41504\,
            in1 => \N__41695\,
            in2 => \N__30905\,
            in3 => \N__25118\,
            lcout => \elapsed_time_ns_1_RNI1BND11_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41696\,
            in1 => \N__25109\,
            in2 => \N__41563\,
            in3 => \N__30629\,
            lcout => \elapsed_time_ns_1_RNIO1ND11_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111111"
        )
    port map (
            in0 => \N__28594\,
            in1 => \N__28580\,
            in2 => \N__28412\,
            in3 => \N__28552\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30841\,
            in2 => \N__25097\,
            in3 => \N__27984\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__25094\,
            in1 => \N__41694\,
            in2 => \N__41549\,
            in3 => \N__30947\,
            lcout => \elapsed_time_ns_1_RNIV8ND11_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_1_c_inv_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28897\,
            in1 => \N__25073\,
            in2 => \N__25085\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_2_c_inv_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25067\,
            in2 => \N__25058\,
            in3 => \N__25487\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_3_c_inv_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25304\,
            in2 => \N__25295\,
            in3 => \N__25460\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_4_c_inv_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25286\,
            in2 => \N__25277\,
            in3 => \N__25442\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_5_c_inv_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25265\,
            in2 => \N__25256\,
            in3 => \N__25658\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_6_c_inv_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25640\,
            in1 => \N__25247\,
            in2 => \N__25238\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_7_c_inv_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25226\,
            in2 => \N__25217\,
            in3 => \N__25622\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_8_c_inv_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25193\,
            in2 => \N__25205\,
            in3 => \N__25604\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_9_c_inv_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25187\,
            in2 => \N__25172\,
            in3 => \N__25586\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_10_c_inv_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25160\,
            in2 => \N__25154\,
            in3 => \N__25568\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_11_c_inv_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25424\,
            in2 => \N__25418\,
            in3 => \N__25550\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_12_c_inv_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25400\,
            in2 => \N__25409\,
            in3 => \N__25532\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_13_c_inv_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25394\,
            in2 => \N__25388\,
            in3 => \N__25811\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_14_c_inv_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25793\,
            in1 => \N__25379\,
            in2 => \N__25373\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_15_c_inv_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25364\,
            in2 => \N__25358\,
            in3 => \N__25775\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_16_c_inv_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25349\,
            in2 => \N__25343\,
            in3 => \N__25754\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_17_c_inv_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25325\,
            in2 => \N__25334\,
            in3 => \N__25736\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_18_c_inv_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25319\,
            in2 => \N__25313\,
            in3 => \N__25718\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_inv_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25514\,
            in2 => \N__25508\,
            in3 => \N__25697\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25499\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNIV5S7_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30800\,
            in2 => \_gnd_net_\,
            in3 => \N__28926\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__28711\,
            in1 => \_gnd_net_\,
            in2 => \N__25496\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJB21_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28712\,
            in2 => \_gnd_net_\,
            in3 => \N__28912\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25493\,
            in2 => \N__28901\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28813\,
            in1 => \N__25486\,
            in2 => \_gnd_net_\,
            in3 => \N__25472\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__45999\,
            ce => 'H',
            sr => \N__45650\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__28822\,
            in1 => \N__25459\,
            in2 => \N__25469\,
            in3 => \N__25445\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__45999\,
            ce => 'H',
            sr => \N__45650\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28814\,
            in1 => \N__25441\,
            in2 => \_gnd_net_\,
            in3 => \N__25427\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__45999\,
            ce => 'H',
            sr => \N__45650\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28823\,
            in1 => \N__25657\,
            in2 => \_gnd_net_\,
            in3 => \N__25643\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__45999\,
            ce => 'H',
            sr => \N__45650\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28815\,
            in1 => \N__25639\,
            in2 => \_gnd_net_\,
            in3 => \N__25625\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__45999\,
            ce => 'H',
            sr => \N__45650\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28824\,
            in1 => \N__25621\,
            in2 => \_gnd_net_\,
            in3 => \N__25607\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__45999\,
            ce => 'H',
            sr => \N__45650\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28816\,
            in1 => \N__25603\,
            in2 => \_gnd_net_\,
            in3 => \N__25589\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__45999\,
            ce => 'H',
            sr => \N__45650\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28870\,
            in1 => \N__25585\,
            in2 => \_gnd_net_\,
            in3 => \N__25571\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_10_25_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__45996\,
            ce => 'H',
            sr => \N__45653\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28817\,
            in1 => \N__25567\,
            in2 => \_gnd_net_\,
            in3 => \N__25553\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__45996\,
            ce => 'H',
            sr => \N__45653\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28867\,
            in1 => \N__25549\,
            in2 => \_gnd_net_\,
            in3 => \N__25535\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__45996\,
            ce => 'H',
            sr => \N__45653\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28818\,
            in1 => \N__25531\,
            in2 => \_gnd_net_\,
            in3 => \N__25517\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__45996\,
            ce => 'H',
            sr => \N__45653\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28868\,
            in1 => \N__25810\,
            in2 => \_gnd_net_\,
            in3 => \N__25796\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__45996\,
            ce => 'H',
            sr => \N__45653\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28819\,
            in1 => \N__25792\,
            in2 => \_gnd_net_\,
            in3 => \N__25778\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__45996\,
            ce => 'H',
            sr => \N__45653\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28869\,
            in1 => \N__25771\,
            in2 => \_gnd_net_\,
            in3 => \N__25757\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__45996\,
            ce => 'H',
            sr => \N__45653\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28820\,
            in1 => \N__25753\,
            in2 => \_gnd_net_\,
            in3 => \N__25739\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__45996\,
            ce => 'H',
            sr => \N__45653\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28866\,
            in1 => \N__25735\,
            in2 => \_gnd_net_\,
            in3 => \N__25721\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_10_26_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__45994\,
            ce => 'H',
            sr => \N__45656\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28828\,
            in1 => \N__25717\,
            in2 => \_gnd_net_\,
            in3 => \N__25703\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__45994\,
            ce => 'H',
            sr => \N__45656\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__25696\,
            in1 => \N__28829\,
            in2 => \_gnd_net_\,
            in3 => \N__25700\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45994\,
            ce => 'H',
            sr => \N__45656\
        );

    \pwm_generator_inst.counter_0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25871\,
            in1 => \N__25681\,
            in2 => \_gnd_net_\,
            in3 => \N__25661\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__46083\,
            ce => 'H',
            sr => \N__45540\
        );

    \pwm_generator_inst.counter_1_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25865\,
            in1 => \N__26074\,
            in2 => \_gnd_net_\,
            in3 => \N__26051\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__46083\,
            ce => 'H',
            sr => \N__45540\
        );

    \pwm_generator_inst.counter_2_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25872\,
            in1 => \N__26047\,
            in2 => \_gnd_net_\,
            in3 => \N__26027\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__46083\,
            ce => 'H',
            sr => \N__45540\
        );

    \pwm_generator_inst.counter_3_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25866\,
            in1 => \N__26020\,
            in2 => \_gnd_net_\,
            in3 => \N__26000\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__46083\,
            ce => 'H',
            sr => \N__45540\
        );

    \pwm_generator_inst.counter_4_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25873\,
            in1 => \N__25996\,
            in2 => \_gnd_net_\,
            in3 => \N__25976\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__46083\,
            ce => 'H',
            sr => \N__45540\
        );

    \pwm_generator_inst.counter_5_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25867\,
            in1 => \N__25971\,
            in2 => \_gnd_net_\,
            in3 => \N__25952\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__46083\,
            ce => 'H',
            sr => \N__45540\
        );

    \pwm_generator_inst.counter_6_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25874\,
            in1 => \N__25948\,
            in2 => \_gnd_net_\,
            in3 => \N__25925\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__46083\,
            ce => 'H',
            sr => \N__45540\
        );

    \pwm_generator_inst.counter_7_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25868\,
            in1 => \N__25921\,
            in2 => \_gnd_net_\,
            in3 => \N__25901\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__46083\,
            ce => 'H',
            sr => \N__45540\
        );

    \pwm_generator_inst.counter_8_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25870\,
            in1 => \N__25897\,
            in2 => \_gnd_net_\,
            in3 => \N__25877\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__46075\,
            ce => 'H',
            sr => \N__45545\
        );

    \pwm_generator_inst.counter_9_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__25831\,
            in1 => \N__25869\,
            in2 => \_gnd_net_\,
            in3 => \N__25835\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46075\,
            ce => 'H',
            sr => \N__45545\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28983\,
            in2 => \_gnd_net_\,
            in3 => \N__28964\,
            lcout => \phase_controller_inst1.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27510\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31294\,
            in2 => \_gnd_net_\,
            in3 => \N__29083\,
            lcout => \phase_controller_inst1.N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36878\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33116\,
            in1 => \N__26134\,
            in2 => \N__26216\,
            in3 => \N__26186\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__27082\,
            in1 => \N__27374\,
            in2 => \N__26162\,
            in3 => \N__27249\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46037\,
            ce => 'H',
            sr => \N__45571\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__27370\,
            in1 => \N__27083\,
            in2 => \N__27256\,
            in3 => \N__26096\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46037\,
            ce => 'H',
            sr => \N__45571\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__27080\,
            in1 => \N__27372\,
            in2 => \N__26087\,
            in3 => \N__27247\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46037\,
            ce => 'H',
            sr => \N__45571\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__27371\,
            in1 => \N__27084\,
            in2 => \N__27257\,
            in3 => \N__26483\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46037\,
            ce => 'H',
            sr => \N__45571\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__27081\,
            in1 => \N__27373\,
            in2 => \N__26474\,
            in3 => \N__27248\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46037\,
            ce => 'H',
            sr => \N__45571\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26460\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26393\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26533\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33112\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26338\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26668\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26272\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26902\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37109\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26804\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26754\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37166\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__26703\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33068\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__26678\,
            in1 => \N__26645\,
            in2 => \N__33125\,
            in3 => \N__26615\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__26594\,
            in1 => \N__26549\,
            in2 => \N__26510\,
            in3 => \N__33069\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__27509\,
            in1 => \N__27586\,
            in2 => \N__33134\,
            in3 => \N__27563\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__27252\,
            in1 => \N__27327\,
            in2 => \N__27119\,
            in3 => \N__27539\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => 'H',
            sr => \N__45588\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__27323\,
            in1 => \N__27254\,
            in2 => \N__27479\,
            in3 => \N__27110\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => 'H',
            sr => \N__45588\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__27250\,
            in1 => \N__27325\,
            in2 => \N__27117\,
            in3 => \N__27470\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => 'H',
            sr => \N__45588\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__27324\,
            in1 => \N__27255\,
            in2 => \N__27419\,
            in3 => \N__27111\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => 'H',
            sr => \N__45588\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__27251\,
            in1 => \N__27326\,
            in2 => \N__27118\,
            in3 => \N__27410\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => 'H',
            sr => \N__45588\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__27322\,
            in1 => \N__27253\,
            in2 => \N__27134\,
            in3 => \N__27109\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => 'H',
            sr => \N__45588\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__28168\,
            in1 => \N__27959\,
            in2 => \N__26891\,
            in3 => \N__27873\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46024\,
            ce => \N__29309\,
            sr => \N__45592\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27871\,
            in1 => \N__28171\,
            in2 => \N__27965\,
            in3 => \N__26863\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46024\,
            ce => \N__29309\,
            sr => \N__45592\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__28169\,
            in1 => \N__27960\,
            in2 => \N__27907\,
            in3 => \N__27874\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46024\,
            ce => \N__29309\,
            sr => \N__45592\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__27872\,
            in1 => \N__28172\,
            in2 => \N__28495\,
            in3 => \N__27760\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46024\,
            ce => \N__29309\,
            sr => \N__45592\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__28167\,
            in1 => \N__27702\,
            in2 => \_gnd_net_\,
            in3 => \N__28313\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46024\,
            ce => \N__29309\,
            sr => \N__45592\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__28311\,
            in1 => \N__28170\,
            in2 => \_gnd_net_\,
            in3 => \N__27677\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46024\,
            ce => \N__29309\,
            sr => \N__45592\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__28066\,
            in1 => \N__28645\,
            in2 => \N__27649\,
            in3 => \N__28312\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46024\,
            ce => \N__29309\,
            sr => \N__45592\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100011101"
        )
    port map (
            in0 => \N__33281\,
            in1 => \N__42191\,
            in2 => \N__33425\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011100"
        )
    port map (
            in0 => \N__33800\,
            in1 => \N__27622\,
            in2 => \N__41564\,
            in3 => \N__30186\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27632\,
            in3 => \N__30281\,
            lcout => \elapsed_time_ns_1_RNIDP2KD1_0_1\,
            ltout => \elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__28056\,
            in1 => \N__27611\,
            in2 => \N__27602\,
            in3 => \N__27598\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46021\,
            ce => \N__29304\,
            sr => \N__45599\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__28308\,
            in1 => \N__28061\,
            in2 => \N__30231\,
            in3 => \N__28166\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46021\,
            ce => \N__29304\,
            sr => \N__45599\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__28163\,
            in1 => \N__41710\,
            in2 => \N__30857\,
            in3 => \N__41530\,
            lcout => \elapsed_time_ns_1_RNIQ4OD11_0_31\,
            ltout => \elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__28306\,
            in1 => \N__28060\,
            in2 => \N__28364\,
            in3 => \N__28354\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46021\,
            ce => \N__29304\,
            sr => \N__45599\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__28164\,
            in1 => \N__28337\,
            in2 => \N__28070\,
            in3 => \N__28309\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46021\,
            ce => \N__29304\,
            sr => \N__45599\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__28307\,
            in1 => \N__28165\,
            in2 => \N__28097\,
            in3 => \N__28062\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46021\,
            ce => \N__29304\,
            sr => \N__45599\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__28019\,
            in1 => \N__41697\,
            in2 => \N__41551\,
            in3 => \N__30881\,
            lcout => \elapsed_time_ns_1_RNIP3OD11_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30856\,
            in1 => \N__45720\,
            in2 => \_gnd_net_\,
            in3 => \N__28006\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__29875\,
            in1 => \N__45718\,
            in2 => \N__27995\,
            in3 => \N__28529\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30471\,
            in1 => \N__30057\,
            in2 => \N__28411\,
            in3 => \N__30336\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__45719\,
            in1 => \N__30855\,
            in2 => \N__28532\,
            in3 => \N__29925\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28378\,
            in2 => \_gnd_net_\,
            in3 => \N__29874\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_382_i\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_382_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__31016\,
            in1 => \N__28520\,
            in2 => \N__28523\,
            in3 => \N__41698\,
            lcout => \elapsed_time_ns_1_RNIS5ND11_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__41699\,
            in1 => \N__28508\,
            in2 => \N__30995\,
            in3 => \N__41511\,
            lcout => \elapsed_time_ns_1_RNIT6ND11_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__28461\,
            in1 => \N__41522\,
            in2 => \N__30305\,
            in3 => \N__41704\,
            lcout => \elapsed_time_ns_1_RNIS4MD11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30684\,
            in1 => \N__30720\,
            in2 => \N__30661\,
            in3 => \N__30750\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__28394\,
            in1 => \N__41703\,
            in2 => \N__41573\,
            in3 => \N__30584\,
            lcout => \elapsed_time_ns_1_RNIQ3ND11_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__45721\,
            in1 => \_gnd_net_\,
            in2 => \N__28382\,
            in3 => \N__29870\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__28643\,
            in1 => \N__41523\,
            in2 => \N__28367\,
            in3 => \N__30122\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__30185\,
            in1 => \_gnd_net_\,
            in2 => \N__28652\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIQURR91_0_3\,
            ltout => \elapsed_time_ns_1_RNIQURR91_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28616\,
            in3 => \N__41386\,
            lcout => \phase_controller_inst1.stoper_hc.N_283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30985\,
            in1 => \N__28538\,
            in2 => \N__31015\,
            in3 => \N__28934\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__30529\,
            in1 => \N__30470\,
            in2 => \_gnd_net_\,
            in3 => \N__30502\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__30301\,
            in1 => \N__28574\,
            in2 => \N__28583\,
            in3 => \N__30335\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30385\,
            in1 => \N__30409\,
            in2 => \N__30439\,
            in3 => \N__30361\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30501\,
            in1 => \N__30528\,
            in2 => \N__28568\,
            in3 => \N__30300\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__30598\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30580\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__30919\,
            in1 => \N__30940\,
            in2 => \_gnd_net_\,
            in3 => \N__30961\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30895\,
            in1 => \N__30622\,
            in2 => \N__30559\,
            in3 => \N__30874\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_2_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__33722\,
            in1 => \N__41830\,
            in2 => \N__41987\,
            in3 => \N__41879\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46000\,
            ce => 'H',
            sr => \N__45639\
        );

    \phase_controller_inst2.stoper_hc.running_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111001001110"
        )
    port map (
            in0 => \N__28713\,
            in1 => \N__28733\,
            in2 => \N__30799\,
            in3 => \N__28927\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46000\,
            ce => 'H',
            sr => \N__45639\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110000001100"
        )
    port map (
            in0 => \N__28928\,
            in1 => \N__41880\,
            in2 => \N__28721\,
            in3 => \N__30795\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46000\,
            ce => 'H',
            sr => \N__45639\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__28821\,
            in1 => \N__28913\,
            in2 => \N__28720\,
            in3 => \N__28896\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46000\,
            ce => 'H',
            sr => \N__45639\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__33747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30791\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__30790\,
            in1 => \N__33746\,
            in2 => \_gnd_net_\,
            in3 => \N__28732\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28691\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46243\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45990\,
            ce => 'H',
            sr => \N__45658\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29018\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43846\,
            in2 => \_gnd_net_\,
            in3 => \N__43925\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29006\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46057\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31238\,
            in2 => \_gnd_net_\,
            in3 => \N__29064\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__28997\,
            in1 => \N__28991\,
            in2 => \N__43678\,
            in3 => \N__43926\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46049\,
            ce => 'H',
            sr => \N__45553\
        );

    \phase_controller_inst1.state_1_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__28985\,
            in1 => \N__31073\,
            in2 => \N__28970\,
            in3 => \N__29104\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46049\,
            ce => 'H',
            sr => \N__45553\
        );

    \phase_controller_inst1.state_2_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__29072\,
            in1 => \N__28969\,
            in2 => \N__31252\,
            in3 => \N__28984\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46049\,
            ce => 'H',
            sr => \N__45553\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__28965\,
            in1 => \N__43897\,
            in2 => \N__43850\,
            in3 => \N__43792\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46043\,
            ce => 'H',
            sr => \N__45558\
        );

    \phase_controller_inst1.start_timer_tr_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__43663\,
            in1 => \N__29050\,
            in2 => \N__32735\,
            in3 => \N__28946\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46043\,
            ce => 'H',
            sr => \N__45558\
        );

    \phase_controller_inst1.state_0_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__29108\,
            in1 => \N__31078\,
            in2 => \N__31298\,
            in3 => \N__29084\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46043\,
            ce => 'H',
            sr => \N__45558\
        );

    \phase_controller_inst1.state_3_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__40517\,
            in1 => \N__29071\,
            in2 => \N__31256\,
            in3 => \N__29051\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46043\,
            ce => 'H',
            sr => \N__45558\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43895\,
            in2 => \_gnd_net_\,
            in3 => \N__29320\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNITEL9_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43845\,
            in2 => \_gnd_net_\,
            in3 => \N__43782\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3D41_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29042\,
            in3 => \N__43896\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3DZ0Z41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__32720\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33245\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29167\,
            in2 => \N__29039\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29273\,
            in1 => \N__29566\,
            in2 => \_gnd_net_\,
            in3 => \N__29030\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__46034\,
            ce => 'H',
            sr => \N__45566\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__29277\,
            in1 => \N__29027\,
            in2 => \N__29537\,
            in3 => \N__29021\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__46034\,
            ce => 'H',
            sr => \N__45566\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29274\,
            in1 => \N__29509\,
            in2 => \_gnd_net_\,
            in3 => \N__29135\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__46034\,
            ce => 'H',
            sr => \N__45566\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29278\,
            in1 => \N__29467\,
            in2 => \_gnd_net_\,
            in3 => \N__29132\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__46034\,
            ce => 'H',
            sr => \N__45566\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29275\,
            in1 => \N__29434\,
            in2 => \_gnd_net_\,
            in3 => \N__29129\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__46034\,
            ce => 'H',
            sr => \N__45566\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29279\,
            in1 => \N__29407\,
            in2 => \_gnd_net_\,
            in3 => \N__29126\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__46034\,
            ce => 'H',
            sr => \N__45566\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29276\,
            in1 => \N__29368\,
            in2 => \_gnd_net_\,
            in3 => \N__29123\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__46034\,
            ce => 'H',
            sr => \N__45566\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29287\,
            in1 => \N__29833\,
            in2 => \_gnd_net_\,
            in3 => \N__29120\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__46032\,
            ce => 'H',
            sr => \N__45572\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29280\,
            in1 => \N__29794\,
            in2 => \_gnd_net_\,
            in3 => \N__29117\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__46032\,
            ce => 'H',
            sr => \N__45572\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29284\,
            in1 => \N__29764\,
            in2 => \_gnd_net_\,
            in3 => \N__29114\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__46032\,
            ce => 'H',
            sr => \N__45572\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29281\,
            in1 => \N__29734\,
            in2 => \_gnd_net_\,
            in3 => \N__29111\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__46032\,
            ce => 'H',
            sr => \N__45572\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29285\,
            in1 => \N__29704\,
            in2 => \_gnd_net_\,
            in3 => \N__29345\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__46032\,
            ce => 'H',
            sr => \N__45572\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29282\,
            in1 => \N__29671\,
            in2 => \_gnd_net_\,
            in3 => \N__29342\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__46032\,
            ce => 'H',
            sr => \N__45572\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29286\,
            in1 => \N__29647\,
            in2 => \_gnd_net_\,
            in3 => \N__29339\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__46032\,
            ce => 'H',
            sr => \N__45572\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29283\,
            in1 => \N__29602\,
            in2 => \_gnd_net_\,
            in3 => \N__29336\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__46032\,
            ce => 'H',
            sr => \N__45572\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29297\,
            in1 => \N__30028\,
            in2 => \_gnd_net_\,
            in3 => \N__29333\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__46028\,
            ce => 'H',
            sr => \N__45577\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29299\,
            in1 => \N__29992\,
            in2 => \_gnd_net_\,
            in3 => \N__29330\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__46028\,
            ce => 'H',
            sr => \N__45577\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29298\,
            in1 => \N__29956\,
            in2 => \_gnd_net_\,
            in3 => \N__29327\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46028\,
            ce => 'H',
            sr => \N__45577\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__43901\,
            in1 => \N__29324\,
            in2 => \N__29168\,
            in3 => \N__29300\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46028\,
            ce => 'H',
            sr => \N__45577\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_1_c_inv_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29183\,
            in2 => \N__29144\,
            in3 => \N__29160\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_2_c_inv_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29579\,
            in2 => \N__29552\,
            in3 => \N__29570\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_3_c_inv_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29543\,
            in2 => \N__29519\,
            in3 => \N__29536\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_4_c_inv_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29510\,
            in1 => \N__29495\,
            in2 => \N__29486\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_5_c_inv_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29477\,
            in2 => \N__29453\,
            in3 => \N__29468\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_6_c_inv_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29444\,
            in2 => \N__29420\,
            in3 => \N__29435\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_7_c_inv_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29408\,
            in1 => \N__29384\,
            in2 => \N__29393\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_8_c_inv_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29354\,
            in2 => \N__29378\,
            in3 => \N__29369\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_9_c_inv_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29846\,
            in2 => \N__29819\,
            in3 => \N__29834\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_10_c_inv_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29780\,
            in2 => \N__29810\,
            in3 => \N__29795\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_11_c_inv_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29750\,
            in2 => \N__29774\,
            in3 => \N__29765\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_12_c_inv_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29720\,
            in2 => \N__29744\,
            in3 => \N__29735\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_13_c_inv_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29690\,
            in2 => \N__29714\,
            in3 => \N__29705\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_14_c_inv_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29684\,
            in2 => \N__29657\,
            in3 => \N__29672\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_15_c_inv_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29648\,
            in1 => \N__29633\,
            in2 => \N__29627\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_16_c_inv_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29615\,
            in2 => \N__29588\,
            in3 => \N__29603\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_17_c_inv_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30041\,
            in2 => \N__30014\,
            in3 => \N__30029\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_18_c_inv_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30005\,
            in2 => \N__29978\,
            in3 => \N__29993\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_inv_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29969\,
            in2 => \N__29942\,
            in3 => \N__29957\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29933\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30121\,
            in1 => \N__33796\,
            in2 => \N__41605\,
            in3 => \N__30131\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30120\,
            in2 => \_gnd_net_\,
            in3 => \N__41601\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__30472\,
            in1 => \N__30130\,
            in2 => \N__29903\,
            in3 => \N__29896\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__30137\,
            in1 => \N__30657\,
            in2 => \N__29879\,
            in3 => \N__30727\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30143\,
            in2 => \_gnd_net_\,
            in3 => \N__30280\,
            lcout => \elapsed_time_ns_1_RNIIU2KD1_0_6\,
            ltout => \elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111010"
        )
    port map (
            in0 => \N__30201\,
            in1 => \N__30059\,
            in2 => \N__30146\,
            in3 => \N__41521\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30058\,
            in1 => \N__30691\,
            in2 => \N__30763\,
            in3 => \N__30340\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30073\,
            in2 => \_gnd_net_\,
            in3 => \N__30097\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31572\,
            in2 => \N__33823\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__46009\,
            ce => \N__33773\,
            sr => \N__45605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31548\,
            in2 => \N__31603\,
            in3 => \N__30086\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__46009\,
            ce => \N__33773\,
            sr => \N__45605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31524\,
            in2 => \N__31577\,
            in3 => \N__30062\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__46009\,
            ce => \N__33773\,
            sr => \N__45605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31815\,
            in2 => \N__31553\,
            in3 => \N__30044\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__46009\,
            ce => \N__33773\,
            sr => \N__45605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31794\,
            in2 => \N__31529\,
            in3 => \N__30515\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__46009\,
            ce => \N__33773\,
            sr => \N__45605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31776\,
            in2 => \N__31820\,
            in3 => \N__30488\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__46009\,
            ce => \N__33773\,
            sr => \N__45605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31795\,
            in2 => \N__31760\,
            in3 => \N__30449\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__46009\,
            ce => \N__33773\,
            sr => \N__45605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31777\,
            in2 => \N__31730\,
            in3 => \N__30422\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__46009\,
            ce => \N__33773\,
            sr => \N__45605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31695\,
            in2 => \N__31759\,
            in3 => \N__30398\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__46003\,
            ce => \N__33771\,
            sr => \N__45619\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31671\,
            in2 => \N__31729\,
            in3 => \N__30374\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__46003\,
            ce => \N__33771\,
            sr => \N__45619\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31647\,
            in2 => \N__31700\,
            in3 => \N__30350\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__46003\,
            ce => \N__33771\,
            sr => \N__45619\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32019\,
            in2 => \N__31676\,
            in3 => \N__30308\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__46003\,
            ce => \N__33771\,
            sr => \N__45619\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31998\,
            in2 => \N__31652\,
            in3 => \N__30284\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__46003\,
            ce => \N__33771\,
            sr => \N__45619\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31980\,
            in2 => \N__32024\,
            in3 => \N__30734\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__46003\,
            ce => \N__33771\,
            sr => \N__45619\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31999\,
            in2 => \N__31964\,
            in3 => \N__30704\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__46003\,
            ce => \N__33771\,
            sr => \N__45619\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31981\,
            in2 => \N__31931\,
            in3 => \N__30668\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__46003\,
            ce => \N__33771\,
            sr => \N__45619\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31901\,
            in2 => \N__31960\,
            in3 => \N__30632\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__45998\,
            ce => \N__33770\,
            sr => \N__45630\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31866\,
            in2 => \N__31930\,
            in3 => \N__30611\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__45998\,
            ce => \N__33770\,
            sr => \N__45630\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31842\,
            in2 => \N__31900\,
            in3 => \N__30587\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__45998\,
            ce => \N__33770\,
            sr => \N__45630\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32346\,
            in2 => \N__31871\,
            in3 => \N__30569\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__45998\,
            ce => \N__33770\,
            sr => \N__45630\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32325\,
            in2 => \N__31847\,
            in3 => \N__30542\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__45998\,
            ce => \N__33770\,
            sr => \N__45630\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32307\,
            in2 => \N__32351\,
            in3 => \N__30998\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__45998\,
            ce => \N__33770\,
            sr => \N__45630\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32326\,
            in2 => \N__32291\,
            in3 => \N__30974\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__45998\,
            ce => \N__33770\,
            sr => \N__45630\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32308\,
            in2 => \N__32261\,
            in3 => \N__30950\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__45998\,
            ce => \N__33770\,
            sr => \N__45630\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32226\,
            in2 => \N__32290\,
            in3 => \N__30929\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_12_23_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__45995\,
            ce => \N__33769\,
            sr => \N__45635\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32202\,
            in2 => \N__32260\,
            in3 => \N__30908\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__45995\,
            ce => \N__33769\,
            sr => \N__45635\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32182\,
            in2 => \N__32231\,
            in3 => \N__30884\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__45995\,
            ce => \N__33769\,
            sr => \N__45635\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32035\,
            in2 => \N__32207\,
            in3 => \N__30863\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__45995\,
            ce => \N__33769\,
            sr => \N__45635\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30860\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45995\,
            ce => \N__33769\,
            sr => \N__45635\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33748\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45993\,
            ce => 'H',
            sr => \N__45640\
        );

    \phase_controller_inst1.S2_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31079\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45991\,
            ce => 'H',
            sr => \N__45651\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45725\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__39895\,
            in1 => \N__32494\,
            in2 => \N__32577\,
            in3 => \N__33997\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46076\,
            ce => \N__44290\,
            sr => \N__45536\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__33995\,
            in1 => \N__39371\,
            in2 => \N__32576\,
            in3 => \N__39896\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46076\,
            ce => \N__44290\,
            sr => \N__45536\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__38592\,
            in1 => \N__32560\,
            in2 => \N__31127\,
            in3 => \N__33996\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46076\,
            ce => \N__44290\,
            sr => \N__45536\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38591\,
            in2 => \_gnd_net_\,
            in3 => \N__35913\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32505\,
            in1 => \N__31103\,
            in2 => \N__39729\,
            in3 => \N__31022\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__31102\,
            in1 => \N__38599\,
            in2 => \N__35924\,
            in3 => \N__32507\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__32506\,
            in1 => \N__39888\,
            in2 => \N__39728\,
            in3 => \N__31101\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111010"
        )
    port map (
            in0 => \N__42737\,
            in1 => \N__39068\,
            in2 => \N__32386\,
            in3 => \N__43168\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31109\,
            in3 => \N__39138\,
            lcout => \elapsed_time_ns_1_RNIUKL2M1_0_6\,
            ltout => \elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__39198\,
            in1 => \N__38966\,
            in2 => \N__31106\,
            in3 => \N__34049\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__39673\,
            in1 => \_gnd_net_\,
            in2 => \N__31091\,
            in3 => \N__34177\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__39889\,
            in1 => \N__32382\,
            in2 => \N__31088\,
            in3 => \N__34001\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46070\,
            ce => \N__44293\,
            sr => \N__45541\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__39919\,
            in1 => \N__43152\,
            in2 => \N__36206\,
            in3 => \N__42741\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__39136\,
            in1 => \_gnd_net_\,
            in2 => \N__31085\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIIJ4DM1_0_19\,
            ltout => \elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39882\,
            in2 => \N__31082\,
            in3 => \N__39731\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46065\,
            ce => \N__44291\,
            sr => \N__45546\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__39730\,
            in1 => \_gnd_net_\,
            in2 => \N__32675\,
            in3 => \N__39886\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46065\,
            ce => \N__44291\,
            sr => \N__45546\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__34223\,
            in1 => \N__39884\,
            in2 => \N__34191\,
            in3 => \N__39732\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46065\,
            ce => \N__44291\,
            sr => \N__45546\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__38976\,
            in1 => \N__39885\,
            in2 => \_gnd_net_\,
            in3 => \N__34000\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46065\,
            ce => \N__44291\,
            sr => \N__45546\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__33998\,
            in1 => \N__39883\,
            in2 => \_gnd_net_\,
            in3 => \N__34051\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46065\,
            ce => \N__44291\,
            sr => \N__45546\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__32362\,
            in1 => \N__33999\,
            in2 => \N__32579\,
            in3 => \N__39887\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46065\,
            ce => \N__44291\,
            sr => \N__45546\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__32764\,
            in1 => \N__32771\,
            in2 => \N__40001\,
            in3 => \N__39734\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46058\,
            ce => \N__39585\,
            sr => \N__45549\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__39873\,
            in1 => \N__39738\,
            in2 => \_gnd_net_\,
            in3 => \N__32823\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46058\,
            ce => \N__39585\,
            sr => \N__45549\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__39739\,
            in1 => \N__39874\,
            in2 => \_gnd_net_\,
            in3 => \N__32674\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46058\,
            ce => \N__39585\,
            sr => \N__45549\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__34007\,
            in1 => \N__31126\,
            in2 => \N__32578\,
            in3 => \N__38603\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46058\,
            ce => \N__39585\,
            sr => \N__45549\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010000"
        )
    port map (
            in0 => \N__32763\,
            in1 => \N__34192\,
            in2 => \N__39200\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33209\,
            in2 => \N__34121\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39587\,
            in1 => \N__34072\,
            in2 => \_gnd_net_\,
            in3 => \N__31154\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__46051\,
            ce => 'H',
            sr => \N__45554\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__39551\,
            in1 => \N__34463\,
            in2 => \N__33167\,
            in3 => \N__31151\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__46051\,
            ce => 'H',
            sr => \N__45554\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39588\,
            in1 => \N__34426\,
            in2 => \_gnd_net_\,
            in3 => \N__31148\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__46051\,
            ce => 'H',
            sr => \N__45554\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39552\,
            in1 => \N__34403\,
            in2 => \_gnd_net_\,
            in3 => \N__31145\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__46051\,
            ce => 'H',
            sr => \N__45554\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39589\,
            in1 => \N__34366\,
            in2 => \_gnd_net_\,
            in3 => \N__31142\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__46051\,
            ce => 'H',
            sr => \N__45554\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39553\,
            in1 => \N__34318\,
            in2 => \_gnd_net_\,
            in3 => \N__31139\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__46051\,
            ce => 'H',
            sr => \N__45554\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39590\,
            in1 => \N__34295\,
            in2 => \_gnd_net_\,
            in3 => \N__31136\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__46051\,
            ce => 'H',
            sr => \N__45554\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39581\,
            in1 => \N__34249\,
            in2 => \_gnd_net_\,
            in3 => \N__31133\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__46045\,
            ce => 'H',
            sr => \N__45559\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39544\,
            in1 => \N__34708\,
            in2 => \_gnd_net_\,
            in3 => \N__31130\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__46045\,
            ce => 'H',
            sr => \N__45559\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39578\,
            in1 => \N__34676\,
            in2 => \_gnd_net_\,
            in3 => \N__31181\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__46045\,
            ce => 'H',
            sr => \N__45559\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39545\,
            in1 => \N__34634\,
            in2 => \_gnd_net_\,
            in3 => \N__31178\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__46045\,
            ce => 'H',
            sr => \N__45559\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39579\,
            in1 => \N__34612\,
            in2 => \_gnd_net_\,
            in3 => \N__31175\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__46045\,
            ce => 'H',
            sr => \N__45559\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39546\,
            in1 => \N__34585\,
            in2 => \_gnd_net_\,
            in3 => \N__31172\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__46045\,
            ce => 'H',
            sr => \N__45559\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39580\,
            in1 => \N__34558\,
            in2 => \_gnd_net_\,
            in3 => \N__31169\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__46045\,
            ce => 'H',
            sr => \N__45559\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39547\,
            in1 => \N__34522\,
            in2 => \_gnd_net_\,
            in3 => \N__31166\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__46045\,
            ce => 'H',
            sr => \N__45559\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39548\,
            in1 => \N__34855\,
            in2 => \_gnd_net_\,
            in3 => \N__31163\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__46038\,
            ce => 'H',
            sr => \N__45562\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39550\,
            in1 => \N__34819\,
            in2 => \_gnd_net_\,
            in3 => \N__31160\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__46038\,
            ce => 'H',
            sr => \N__45562\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39549\,
            in1 => \N__34798\,
            in2 => \_gnd_net_\,
            in3 => \N__31157\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46038\,
            ce => 'H',
            sr => \N__45562\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101011001010"
        )
    port map (
            in0 => \N__31287\,
            in1 => \N__33244\,
            in2 => \N__33203\,
            in3 => \N__34772\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46038\,
            ce => 'H',
            sr => \N__45562\
        );

    \phase_controller_inst2.state_0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__43740\,
            in1 => \N__31270\,
            in2 => \N__46247\,
            in3 => \N__46152\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46035\,
            ce => 'H',
            sr => \N__45567\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__31271\,
            in1 => \N__43508\,
            in2 => \N__43583\,
            in3 => \N__43616\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46035\,
            ce => 'H',
            sr => \N__45567\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31269\,
            in2 => \_gnd_net_\,
            in3 => \N__46151\,
            lcout => \phase_controller_inst2.time_passed_RNI9M3O\,
            ltout => \phase_controller_inst2.time_passed_RNI9M3O_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_3_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__41946\,
            in1 => \N__40513\,
            in2 => \N__31259\,
            in3 => \N__33715\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46035\,
            ce => 'H',
            sr => \N__45567\
        );

    \phase_controller_inst1.state_4_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__40564\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43650\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46035\,
            ce => 'H',
            sr => \N__45567\
        );

    \current_shift_inst.stop_timer_s1_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__31253\,
            in1 => \N__31195\,
            in2 => \N__31507\,
            in3 => \N__32423\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46033\,
            ce => 'H',
            sr => \N__45573\
        );

    \current_shift_inst.timer_s1.running_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__31502\,
            in1 => \N__35810\,
            in2 => \_gnd_net_\,
            in3 => \N__32424\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46033\,
            ce => 'H',
            sr => \N__45573\
        );

    \current_shift_inst.start_timer_s1_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__31194\,
            in1 => \N__31503\,
            in2 => \_gnd_net_\,
            in3 => \N__31255\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46033\,
            ce => 'H',
            sr => \N__45573\
        );

    \phase_controller_inst1.S1_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31254\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46033\,
            ce => 'H',
            sr => \N__45573\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31448\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31401\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31334\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33263\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37565\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46030\,
            ce => \N__41021\,
            sr => \N__45578\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35381\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35336\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__47194\,
            in1 => \N__33385\,
            in2 => \N__44054\,
            in3 => \N__31480\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37532\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46025\,
            ce => \N__41020\,
            sr => \N__45582\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31475\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__33386\,
            in1 => \N__47195\,
            in2 => \N__31481\,
            in3 => \N__44053\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__42192\,
            in1 => \N__33384\,
            in2 => \_gnd_net_\,
            in3 => \N__31476\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47196\,
            in2 => \_gnd_net_\,
            in3 => \N__33553\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__47197\,
            in1 => \_gnd_net_\,
            in2 => \N__33557\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42241\,
            in1 => \N__36768\,
            in2 => \_gnd_net_\,
            in3 => \N__36726\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46975\,
            in1 => \N__47325\,
            in2 => \N__35344\,
            in3 => \N__33310\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42239\,
            in1 => \N__35382\,
            in2 => \_gnd_net_\,
            in3 => \N__33339\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__46973\,
            in1 => \N__47327\,
            in2 => \N__35200\,
            in3 => \N__35473\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__42238\,
            in1 => \N__33367\,
            in2 => \_gnd_net_\,
            in3 => \N__35436\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35337\,
            in1 => \N__42240\,
            in2 => \_gnd_net_\,
            in3 => \N__33309\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__47326\,
            in1 => \N__46976\,
            in2 => \N__36773\,
            in3 => \N__36727\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__46974\,
            in1 => \N__47328\,
            in2 => \N__35201\,
            in3 => \N__35474\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44917\,
            in1 => \N__47335\,
            in2 => \N__47003\,
            in3 => \N__44878\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__31508\,
            in1 => \N__35817\,
            in2 => \_gnd_net_\,
            in3 => \N__32428\,
            lcout => \current_shift_inst.timer_s1.N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44916\,
            in1 => \N__47334\,
            in2 => \_gnd_net_\,
            in3 => \N__44877\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__47333\,
            in1 => \N__46992\,
            in2 => \N__47450\,
            in3 => \N__47470\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44915\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47332\,
            in1 => \N__41340\,
            in2 => \_gnd_net_\,
            in3 => \N__41292\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45228\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__36981\,
            in1 => \N__42257\,
            in2 => \_gnd_net_\,
            in3 => \N__42387\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37061\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35278\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45075\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47336\,
            in1 => \N__44680\,
            in2 => \N__47004\,
            in3 => \N__44698\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32143\,
            in1 => \N__33816\,
            in2 => \_gnd_net_\,
            in3 => \N__31613\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__46010\,
            ce => \N__32471\,
            sr => \N__45606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32139\,
            in1 => \N__31596\,
            in2 => \_gnd_net_\,
            in3 => \N__31580\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__46010\,
            ce => \N__32471\,
            sr => \N__45606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32144\,
            in1 => \N__31573\,
            in2 => \_gnd_net_\,
            in3 => \N__31556\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__46010\,
            ce => \N__32471\,
            sr => \N__45606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32140\,
            in1 => \N__31549\,
            in2 => \_gnd_net_\,
            in3 => \N__31532\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__46010\,
            ce => \N__32471\,
            sr => \N__45606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32145\,
            in1 => \N__31525\,
            in2 => \_gnd_net_\,
            in3 => \N__31823\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__46010\,
            ce => \N__32471\,
            sr => \N__45606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32141\,
            in1 => \N__31816\,
            in2 => \_gnd_net_\,
            in3 => \N__31799\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__46010\,
            ce => \N__32471\,
            sr => \N__45606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32146\,
            in1 => \N__31796\,
            in2 => \_gnd_net_\,
            in3 => \N__31781\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__46010\,
            ce => \N__32471\,
            sr => \N__45606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32142\,
            in1 => \N__31778\,
            in2 => \_gnd_net_\,
            in3 => \N__31763\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__46010\,
            ce => \N__32471\,
            sr => \N__45606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32150\,
            in1 => \N__31752\,
            in2 => \_gnd_net_\,
            in3 => \N__31733\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__46004\,
            ce => \N__32469\,
            sr => \N__45620\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32162\,
            in1 => \N__31722\,
            in2 => \_gnd_net_\,
            in3 => \N__31703\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__46004\,
            ce => \N__32469\,
            sr => \N__45620\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32147\,
            in1 => \N__31696\,
            in2 => \_gnd_net_\,
            in3 => \N__31679\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__46004\,
            ce => \N__32469\,
            sr => \N__45620\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32159\,
            in1 => \N__31672\,
            in2 => \_gnd_net_\,
            in3 => \N__31655\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__46004\,
            ce => \N__32469\,
            sr => \N__45620\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32148\,
            in1 => \N__31648\,
            in2 => \_gnd_net_\,
            in3 => \N__31631\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__46004\,
            ce => \N__32469\,
            sr => \N__45620\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32160\,
            in1 => \N__32020\,
            in2 => \_gnd_net_\,
            in3 => \N__32003\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__46004\,
            ce => \N__32469\,
            sr => \N__45620\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32149\,
            in1 => \N__32000\,
            in2 => \_gnd_net_\,
            in3 => \N__31985\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__46004\,
            ce => \N__32469\,
            sr => \N__45620\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32161\,
            in1 => \N__31982\,
            in2 => \_gnd_net_\,
            in3 => \N__31967\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__46004\,
            ce => \N__32469\,
            sr => \N__45620\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32155\,
            in1 => \N__31953\,
            in2 => \_gnd_net_\,
            in3 => \N__31934\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__46001\,
            ce => \N__32470\,
            sr => \N__45631\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32165\,
            in1 => \N__31923\,
            in2 => \_gnd_net_\,
            in3 => \N__31904\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__46001\,
            ce => \N__32470\,
            sr => \N__45631\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32156\,
            in1 => \N__31893\,
            in2 => \_gnd_net_\,
            in3 => \N__31874\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__46001\,
            ce => \N__32470\,
            sr => \N__45631\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32166\,
            in1 => \N__31867\,
            in2 => \_gnd_net_\,
            in3 => \N__31850\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__46001\,
            ce => \N__32470\,
            sr => \N__45631\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32157\,
            in1 => \N__31843\,
            in2 => \_gnd_net_\,
            in3 => \N__31826\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__46001\,
            ce => \N__32470\,
            sr => \N__45631\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32167\,
            in1 => \N__32347\,
            in2 => \_gnd_net_\,
            in3 => \N__32330\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__46001\,
            ce => \N__32470\,
            sr => \N__45631\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32158\,
            in1 => \N__32327\,
            in2 => \_gnd_net_\,
            in3 => \N__32312\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__46001\,
            ce => \N__32470\,
            sr => \N__45631\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32168\,
            in1 => \N__32309\,
            in2 => \_gnd_net_\,
            in3 => \N__32294\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__46001\,
            ce => \N__32470\,
            sr => \N__45631\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32151\,
            in1 => \N__32283\,
            in2 => \_gnd_net_\,
            in3 => \N__32264\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__45997\,
            ce => \N__32462\,
            sr => \N__45636\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32163\,
            in1 => \N__32253\,
            in2 => \_gnd_net_\,
            in3 => \N__32234\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__45997\,
            ce => \N__32462\,
            sr => \N__45636\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32152\,
            in1 => \N__32227\,
            in2 => \_gnd_net_\,
            in3 => \N__32210\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__45997\,
            ce => \N__32462\,
            sr => \N__45636\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32164\,
            in1 => \N__32203\,
            in2 => \_gnd_net_\,
            in3 => \N__32186\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__45997\,
            ce => \N__32462\,
            sr => \N__45636\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32153\,
            in1 => \N__32183\,
            in2 => \_gnd_net_\,
            in3 => \N__32171\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__45997\,
            ce => \N__32462\,
            sr => \N__45636\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__32036\,
            in1 => \N__32154\,
            in2 => \_gnd_net_\,
            in3 => \N__32039\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45997\,
            ce => \N__32462\,
            sr => \N__45636\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35818\,
            in2 => \_gnd_net_\,
            in3 => \N__32429\,
            lcout => \current_shift_inst.timer_s1.N_166_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111011111110"
        )
    port map (
            in0 => \N__42733\,
            in1 => \N__32610\,
            in2 => \N__43172\,
            in3 => \N__38657\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32393\,
            in3 => \N__39133\,
            lcout => \elapsed_time_ns_1_RNIPFL2M1_0_1\,
            ltout => \elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__32551\,
            in1 => \N__32596\,
            in2 => \N__32390\,
            in3 => \N__32618\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46084\,
            ce => \N__39598\,
            sr => \N__45531\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__33992\,
            in1 => \N__39894\,
            in2 => \N__32387\,
            in3 => \N__32559\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46084\,
            ce => \N__39598\,
            sr => \N__45531\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__39891\,
            in1 => \N__32363\,
            in2 => \N__32574\,
            in3 => \N__33993\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46084\,
            ce => \N__39598\,
            sr => \N__45531\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__33991\,
            in1 => \N__39893\,
            in2 => \N__32495\,
            in3 => \N__32558\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46084\,
            ce => \N__39598\,
            sr => \N__45531\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__39892\,
            in1 => \N__39370\,
            in2 => \N__32575\,
            in3 => \N__33994\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46084\,
            ce => \N__39598\,
            sr => \N__45531\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111000"
        )
    port map (
            in0 => \N__39017\,
            in1 => \N__43156\,
            in2 => \N__42745\,
            in3 => \N__32753\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__42824\,
            in1 => \N__42971\,
            in2 => \N__43169\,
            in3 => \N__34169\,
            lcout => \elapsed_time_ns_1_RNIUCHF91_0_15\,
            ltout => \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40080\,
            in2 => \N__32636\,
            in3 => \N__32754\,
            lcout => \phase_controller_inst1.stoper_tr.N_251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32633\,
            in2 => \_gnd_net_\,
            in3 => \N__39137\,
            lcout => \elapsed_time_ns_1_RNI1OL2M1_0_9\,
            ltout => \elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40081\,
            in2 => \N__32627\,
            in3 => \N__39199\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.N_211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__34220\,
            in1 => \N__34170\,
            in2 => \N__32624\,
            in3 => \N__39677\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32611\,
            in2 => \N__32621\,
            in3 => \N__39890\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__32612\,
            in1 => \N__32597\,
            in2 => \N__32582\,
            in3 => \N__32567\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46077\,
            ce => \N__44294\,
            sr => \N__45537\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32684\,
            in1 => \N__39918\,
            in2 => \N__32795\,
            in3 => \N__34026\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__43146\,
            in1 => \N__32484\,
            in2 => \N__42994\,
            in3 => \N__35867\,
            lcout => \elapsed_time_ns_1_RNICG2591_0_4\,
            ltout => \elapsed_time_ns_1_RNICG2591_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32668\,
            in1 => \N__32822\,
            in2 => \N__32687\,
            in3 => \N__39356\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__43148\,
            in1 => \N__36365\,
            in2 => \N__42746\,
            in3 => \N__32670\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__39135\,
            in1 => \_gnd_net_\,
            in2 => \N__32678\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIFG4DM1_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32645\,
            in2 => \_gnd_net_\,
            in3 => \N__39134\,
            lcout => \elapsed_time_ns_1_RNIGH4DM1_0_17\,
            ltout => \elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__32669\,
            in1 => \N__39917\,
            in2 => \N__32648\,
            in3 => \N__34025\,
            lcout => \phase_controller_inst1.stoper_tr.N_214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__43147\,
            in1 => \N__34052\,
            in2 => \N__42995\,
            in3 => \N__39044\,
            lcout => \elapsed_time_ns_1_RNIGK2591_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__36316\,
            in1 => \N__42735\,
            in2 => \N__32830\,
            in3 => \N__43157\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__42736\,
            in1 => \N__34027\,
            in2 => \N__43171\,
            in3 => \N__36257\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39140\,
            in2 => \N__32639\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIHI4DM1_0_18\,
            ltout => \elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__39736\,
            in1 => \_gnd_net_\,
            in2 => \N__32834\,
            in3 => \N__39860\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46066\,
            ce => \N__44289\,
            sr => \N__45547\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__39859\,
            in1 => \_gnd_net_\,
            in2 => \N__32831\,
            in3 => \N__39737\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46066\,
            ce => \N__44289\,
            sr => \N__45547\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__43430\,
            in1 => \N__42990\,
            in2 => \N__43170\,
            in3 => \N__39858\,
            lcout => \elapsed_time_ns_1_RNISCJF91_0_31\,
            ltout => \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111110"
        )
    port map (
            in0 => \N__32801\,
            in1 => \N__32794\,
            in2 => \N__32774\,
            in3 => \N__39735\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__32765\,
            in1 => \N__39733\,
            in2 => \N__32738\,
            in3 => \N__39993\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46066\,
            ce => \N__44289\,
            sr => \N__45547\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32730\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46059\,
            ce => 'H',
            sr => \N__45550\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__33199\,
            in1 => \N__33179\,
            in2 => \N__34120\,
            in3 => \N__39586\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46059\,
            ce => 'H',
            sr => \N__45550\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__33232\,
            in1 => \N__32695\,
            in2 => \_gnd_net_\,
            in3 => \N__32734\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => \phase_controller_inst1.stoper_tr.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101011111010"
        )
    port map (
            in0 => \N__32696\,
            in1 => \N__34771\,
            in2 => \N__32699\,
            in3 => \N__33234\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46052\,
            ce => 'H',
            sr => \N__45555\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIJPMR_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__33233\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34767\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33212\,
            in3 => \N__33197\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6N32_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33198\,
            in2 => \_gnd_net_\,
            in3 => \N__33178\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6NZ0Z32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46613\,
            in1 => \N__47180\,
            in2 => \N__41353\,
            in3 => \N__41302\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__47177\,
            in1 => \N__42395\,
            in2 => \N__36986\,
            in3 => \N__46617\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46618\,
            in1 => \N__47178\,
            in2 => \N__35294\,
            in3 => \N__35245\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37079\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35519\,
            in1 => \N__47179\,
            in2 => \N__46802\,
            in3 => \N__35135\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33143\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47046\,
            in1 => \N__47109\,
            in2 => \_gnd_net_\,
            in3 => \N__46389\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41053\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46039\,
            ce => \N__41022\,
            sr => \N__45563\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46605\,
            in1 => \N__47105\,
            in2 => \N__35441\,
            in3 => \N__33373\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100011"
        )
    port map (
            in0 => \N__33374\,
            in1 => \N__35437\,
            in2 => \N__47193\,
            in3 => \N__46606\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__33277\,
            in1 => \N__33290\,
            in2 => \_gnd_net_\,
            in3 => \N__47104\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33421\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47103\,
            in2 => \N__33284\,
            in3 => \N__33276\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45080\,
            in1 => \N__47204\,
            in2 => \N__46806\,
            in3 => \N__45036\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47198\,
            in1 => \N__42044\,
            in2 => \N__46805\,
            in3 => \N__42010\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46632\,
            in1 => \N__47199\,
            in2 => \N__35399\,
            in3 => \N__33344\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47205\,
            in1 => \N__35515\,
            in2 => \N__46804\,
            in3 => \N__35134\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46633\,
            in1 => \N__47200\,
            in2 => \N__35348\,
            in3 => \N__33314\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__47203\,
            in1 => \N__46628\,
            in2 => \N__42445\,
            in3 => \N__42487\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__35246\,
            in1 => \N__47201\,
            in2 => \N__46807\,
            in3 => \N__35293\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47202\,
            in1 => \N__35572\,
            in2 => \N__46803\,
            in3 => \N__35114\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__47223\,
            in1 => \N__46879\,
            in2 => \N__35573\,
            in3 => \N__35113\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__46881\,
            in1 => \N__47225\,
            in2 => \N__41749\,
            in3 => \N__41785\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__47226\,
            in1 => \N__46882\,
            in2 => \N__45239\,
            in3 => \N__45190\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46883\,
            in1 => \N__47227\,
            in2 => \N__41231\,
            in3 => \N__41261\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__47222\,
            in1 => \N__46885\,
            in2 => \N__42081\,
            in3 => \N__42121\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46880\,
            in1 => \N__47224\,
            in2 => \N__45154\,
            in3 => \N__45112\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__47221\,
            in1 => \N__46884\,
            in2 => \N__35395\,
            in3 => \N__33340\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46878\,
            in1 => \N__47228\,
            in2 => \N__42341\,
            in3 => \N__42292\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33431\,
            in2 => \N__33417\,
            in3 => \N__33410\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35150\,
            in2 => \_gnd_net_\,
            in3 => \N__33356\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35252\,
            in2 => \_gnd_net_\,
            in3 => \N__33353\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33350\,
            in2 => \_gnd_net_\,
            in3 => \N__33323\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33320\,
            in2 => \_gnd_net_\,
            in3 => \N__33296\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35210\,
            in2 => \_gnd_net_\,
            in3 => \N__33293\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42353\,
            in2 => \_gnd_net_\,
            in3 => \N__33482\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33542\,
            in2 => \_gnd_net_\,
            in3 => \N__33479\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33476\,
            in2 => \_gnd_net_\,
            in3 => \N__33461\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33632\,
            in2 => \_gnd_net_\,
            in3 => \N__33458\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33653\,
            in2 => \_gnd_net_\,
            in3 => \N__33455\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33527\,
            in2 => \_gnd_net_\,
            in3 => \N__33452\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33449\,
            in2 => \_gnd_net_\,
            in3 => \N__33440\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33608\,
            in2 => \_gnd_net_\,
            in3 => \N__33437\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33641\,
            in2 => \_gnd_net_\,
            in3 => \N__33434\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33518\,
            in2 => \_gnd_net_\,
            in3 => \N__33509\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33533\,
            in2 => \_gnd_net_\,
            in3 => \N__33506\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33617\,
            in2 => \_gnd_net_\,
            in3 => \N__33503\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33662\,
            in2 => \_gnd_net_\,
            in3 => \N__33500\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33599\,
            in2 => \_gnd_net_\,
            in3 => \N__33497\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33590\,
            in2 => \_gnd_net_\,
            in3 => \N__33494\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37577\,
            in2 => \_gnd_net_\,
            in3 => \N__33491\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33860\,
            in2 => \_gnd_net_\,
            in3 => \N__33488\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33842\,
            in2 => \_gnd_net_\,
            in3 => \N__33485\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33623\,
            in2 => \_gnd_net_\,
            in3 => \N__33581\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33851\,
            in2 => \_gnd_net_\,
            in3 => \N__33578\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33833\,
            in2 => \_gnd_net_\,
            in3 => \N__33575\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35837\,
            in2 => \_gnd_net_\,
            in3 => \N__33572\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33569\,
            in2 => \_gnd_net_\,
            in3 => \N__33563\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33560\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42101\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41211\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42467\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47429\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45131\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35499\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35550\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44978\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35457\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41768\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44663\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41101\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44756\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41321\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44840\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47027\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33824\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46005\,
            ce => \N__33772\,
            sr => \N__45621\
        );

    \phase_controller_inst2.start_timer_hc_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__43677\,
            in1 => \N__35825\,
            in2 => \N__33749\,
            in3 => \N__33683\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46002\,
            ce => 'H',
            sr => \N__45632\
        );

    \phase_controller_inst2.start_timer_hc_RNO_1_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41962\,
            in2 => \_gnd_net_\,
            in3 => \N__33714\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35741\,
            in2 => \_gnd_net_\,
            in3 => \N__46355\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_434_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35696\,
            in1 => \N__38715\,
            in2 => \_gnd_net_\,
            in3 => \N__33665\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_5_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__46102\,
            ce => \N__35785\,
            sr => \N__45519\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35683\,
            in1 => \N__35886\,
            in2 => \_gnd_net_\,
            in3 => \N__33887\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__46102\,
            ce => \N__35785\,
            sr => \N__45519\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35697\,
            in1 => \N__36144\,
            in2 => \_gnd_net_\,
            in3 => \N__33884\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__46102\,
            ce => \N__35785\,
            sr => \N__45519\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35684\,
            in1 => \N__36123\,
            in2 => \_gnd_net_\,
            in3 => \N__33881\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__46102\,
            ce => \N__35785\,
            sr => \N__45519\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35698\,
            in1 => \N__36099\,
            in2 => \_gnd_net_\,
            in3 => \N__33878\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__46102\,
            ce => \N__35785\,
            sr => \N__45519\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35685\,
            in1 => \N__36072\,
            in2 => \_gnd_net_\,
            in3 => \N__33875\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__46102\,
            ce => \N__35785\,
            sr => \N__45519\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35699\,
            in1 => \N__36042\,
            in2 => \_gnd_net_\,
            in3 => \N__33872\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__46102\,
            ce => \N__35785\,
            sr => \N__45519\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35686\,
            in1 => \N__36015\,
            in2 => \_gnd_net_\,
            in3 => \N__33869\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__46102\,
            ce => \N__35785\,
            sr => \N__45519\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35717\,
            in1 => \N__35988\,
            in2 => \_gnd_net_\,
            in3 => \N__33866\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_6_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__46097\,
            ce => \N__35777\,
            sr => \N__45526\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35674\,
            in1 => \N__35955\,
            in2 => \_gnd_net_\,
            in3 => \N__33863\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__46097\,
            ce => \N__35777\,
            sr => \N__45526\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35714\,
            in1 => \N__36456\,
            in2 => \_gnd_net_\,
            in3 => \N__33914\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__46097\,
            ce => \N__35777\,
            sr => \N__45526\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35671\,
            in1 => \N__36432\,
            in2 => \_gnd_net_\,
            in3 => \N__33911\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__46097\,
            ce => \N__35777\,
            sr => \N__45526\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35715\,
            in1 => \N__36405\,
            in2 => \_gnd_net_\,
            in3 => \N__33908\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__46097\,
            ce => \N__35777\,
            sr => \N__45526\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35672\,
            in1 => \N__36381\,
            in2 => \_gnd_net_\,
            in3 => \N__33905\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__46097\,
            ce => \N__35777\,
            sr => \N__45526\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35716\,
            in1 => \N__36333\,
            in2 => \_gnd_net_\,
            in3 => \N__33902\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__46097\,
            ce => \N__35777\,
            sr => \N__45526\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35673\,
            in1 => \N__36271\,
            in2 => \_gnd_net_\,
            in3 => \N__33899\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__46097\,
            ce => \N__35777\,
            sr => \N__45526\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35675\,
            in1 => \N__36225\,
            in2 => \_gnd_net_\,
            in3 => \N__33896\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__46092\,
            ce => \N__35786\,
            sr => \N__45528\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35679\,
            in1 => \N__36168\,
            in2 => \_gnd_net_\,
            in3 => \N__33893\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__46092\,
            ce => \N__35786\,
            sr => \N__45528\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35676\,
            in1 => \N__36711\,
            in2 => \_gnd_net_\,
            in3 => \N__33890\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__46092\,
            ce => \N__35786\,
            sr => \N__45528\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35680\,
            in1 => \N__36690\,
            in2 => \_gnd_net_\,
            in3 => \N__33941\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__46092\,
            ce => \N__35786\,
            sr => \N__45528\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35677\,
            in1 => \N__36666\,
            in2 => \_gnd_net_\,
            in3 => \N__33938\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__46092\,
            ce => \N__35786\,
            sr => \N__45528\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35681\,
            in1 => \N__36639\,
            in2 => \_gnd_net_\,
            in3 => \N__33935\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__46092\,
            ce => \N__35786\,
            sr => \N__45528\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35678\,
            in1 => \N__36609\,
            in2 => \_gnd_net_\,
            in3 => \N__33932\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__46092\,
            ce => \N__35786\,
            sr => \N__45528\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35682\,
            in1 => \N__36582\,
            in2 => \_gnd_net_\,
            in3 => \N__33929\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__46092\,
            ce => \N__35786\,
            sr => \N__45528\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35718\,
            in1 => \N__36555\,
            in2 => \_gnd_net_\,
            in3 => \N__33926\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__46085\,
            ce => \N__35784\,
            sr => \N__45532\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35722\,
            in1 => \N__36522\,
            in2 => \_gnd_net_\,
            in3 => \N__33923\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__46085\,
            ce => \N__35784\,
            sr => \N__45532\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35719\,
            in1 => \N__36498\,
            in2 => \_gnd_net_\,
            in3 => \N__33920\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__46085\,
            ce => \N__35784\,
            sr => \N__45532\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35723\,
            in1 => \N__36834\,
            in2 => \_gnd_net_\,
            in3 => \N__33917\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__46085\,
            ce => \N__35784\,
            sr => \N__45532\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35720\,
            in1 => \N__36475\,
            in2 => \_gnd_net_\,
            in3 => \N__34058\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__46085\,
            ce => \N__35784\,
            sr => \N__45532\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__36853\,
            in1 => \N__35721\,
            in2 => \_gnd_net_\,
            in3 => \N__34055\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46085\,
            ce => \N__35784\,
            sr => \N__45532\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__39876\,
            in1 => \N__34050\,
            in2 => \_gnd_net_\,
            in3 => \N__34003\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46078\,
            ce => \N__39599\,
            sr => \N__45538\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__34028\,
            in1 => \N__39879\,
            in2 => \_gnd_net_\,
            in3 => \N__39751\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46078\,
            ce => \N__39599\,
            sr => \N__45538\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__39875\,
            in1 => \N__38977\,
            in2 => \_gnd_net_\,
            in3 => \N__34002\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46078\,
            ce => \N__39599\,
            sr => \N__45538\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__39990\,
            in1 => \N__39880\,
            in2 => \N__39236\,
            in3 => \N__39752\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46078\,
            ce => \N__39599\,
            sr => \N__45538\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__39877\,
            in1 => \N__39991\,
            in2 => \N__39754\,
            in3 => \N__43336\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46078\,
            ce => \N__39599\,
            sr => \N__45538\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__39878\,
            in1 => \N__39992\,
            in2 => \N__39755\,
            in3 => \N__39262\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46078\,
            ce => \N__39599\,
            sr => \N__45538\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__34222\,
            in1 => \N__39881\,
            in2 => \N__34190\,
            in3 => \N__39753\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46078\,
            ce => \N__39599\,
            sr => \N__45538\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__39863\,
            in1 => \N__40076\,
            in2 => \N__40000\,
            in3 => \N__39744\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46071\,
            ce => \N__44292\,
            sr => \N__45542\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__40075\,
            in1 => \N__43167\,
            in2 => \N__42789\,
            in3 => \N__42734\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34226\,
            in3 => \N__39139\,
            lcout => \elapsed_time_ns_1_RNIDE4DM1_0_14\,
            ltout => \elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34221\,
            in2 => \N__34199\,
            in3 => \N__34196\,
            lcout => \phase_controller_inst1.stoper_tr.N_241\,
            ltout => \phase_controller_inst1.stoper_tr.N_241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__39861\,
            in1 => \N__43337\,
            in2 => \N__34136\,
            in3 => \N__39742\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46071\,
            ce => \N__44292\,
            sr => \N__45542\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__39740\,
            in1 => \N__39864\,
            in2 => \N__39266\,
            in3 => \N__39988\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46071\,
            ce => \N__44292\,
            sr => \N__45542\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__39862\,
            in1 => \N__39232\,
            in2 => \N__39999\,
            in3 => \N__39743\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46071\,
            ce => \N__44292\,
            sr => \N__45542\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__39741\,
            in1 => \N__39865\,
            in2 => \N__40028\,
            in3 => \N__39989\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46071\,
            ce => \N__44292\,
            sr => \N__45542\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_1_c_inv_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34133\,
            in2 => \N__34094\,
            in3 => \N__34110\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_2_c_inv_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34085\,
            in2 => \N__34487\,
            in3 => \N__34073\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_3_c_inv_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34475\,
            in2 => \N__34448\,
            in3 => \N__34462\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_4_c_inv_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34439\,
            in2 => \N__34412\,
            in3 => \N__34427\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_5_c_inv_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34402\,
            in1 => \N__34388\,
            in2 => \N__34376\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_6_c_inv_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34367\,
            in1 => \N__34352\,
            in2 => \N__34340\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_7_c_inv_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34328\,
            in2 => \N__34304\,
            in3 => \N__34319\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_8_c_inv_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34294\,
            in1 => \N__34280\,
            in2 => \N__34271\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_9_c_inv_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34262\,
            in2 => \N__34235\,
            in3 => \N__34250\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_10_c_inv_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34718\,
            in2 => \N__34694\,
            in3 => \N__34709\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_11_c_inv_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34685\,
            in2 => \N__34661\,
            in3 => \N__34675\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_12_c_inv_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34619\,
            in2 => \N__34649\,
            in3 => \N__34633\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_13_c_inv_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34613\,
            in1 => \N__39938\,
            in2 => \N__34598\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_14_c_inv_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34586\,
            in1 => \N__40052\,
            in2 => \N__34571\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_15_c_inv_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34559\,
            in1 => \N__34544\,
            in2 => \N__34532\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_16_c_inv_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34523\,
            in1 => \N__34508\,
            in2 => \N__34496\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_17_c_inv_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34868\,
            in2 => \N__34841\,
            in3 => \N__34856\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_18_c_inv_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34805\,
            in2 => \N__34832\,
            in3 => \N__34820\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_inv_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39611\,
            in2 => \N__34784\,
            in3 => \N__34799\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34775\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__43573\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43529\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34751\,
            in2 => \N__44095\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44040\,
            in2 => \N__34745\,
            in3 => \N__37215\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37216\,
            in1 => \N__46509\,
            in2 => \N__34730\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34940\,
            in2 => \N__46648\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46513\,
            in2 => \N__34934\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34925\,
            in2 => \N__46649\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46517\,
            in2 => \N__34919\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34904\,
            in2 => \N__46650\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46554\,
            in2 => \N__34898\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34889\,
            in2 => \N__46756\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46558\,
            in2 => \N__34883\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34874\,
            in2 => \N__46757\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46562\,
            in2 => \N__35012\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35003\,
            in2 => \N__46758\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46566\,
            in2 => \N__34997\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34988\,
            in2 => \N__46759\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46760\,
            in2 => \N__34982\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34973\,
            in2 => \N__46911\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46764\,
            in2 => \N__34967\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34952\,
            in2 => \N__46912\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46768\,
            in2 => \N__35090\,
            in3 => \N__35075\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41129\,
            in2 => \N__46913\,
            in3 => \N__35072\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46772\,
            in2 => \N__35069\,
            in3 => \N__35060\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35219\,
            in2 => \N__46914\,
            in3 => \N__35057\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46776\,
            in2 => \N__35144\,
            in3 => \N__35054\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35180\,
            in2 => \N__46915\,
            in3 => \N__35051\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46780\,
            in2 => \N__35048\,
            in3 => \N__35033\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35030\,
            in2 => \N__46916\,
            in3 => \N__35018\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46784\,
            in2 => \N__40757\,
            in3 => \N__35015\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35171\,
            in2 => \N__46917\,
            in3 => \N__35159\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46788\,
            in2 => \N__44539\,
            in3 => \N__35156\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_0_11_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110100100111"
        )
    port map (
            in0 => \N__40937\,
            in1 => \N__41138\,
            in2 => \N__44498\,
            in3 => \N__35153\,
            lcout => \current_shift_inst.control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35427\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41778\,
            in1 => \N__42248\,
            in2 => \_gnd_net_\,
            in3 => \N__41733\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__47352\,
            in1 => \N__46886\,
            in2 => \N__44857\,
            in3 => \N__44811\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42039\,
            in1 => \N__42245\,
            in2 => \_gnd_net_\,
            in3 => \N__42003\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42249\,
            in1 => \N__35508\,
            in2 => \_gnd_net_\,
            in3 => \N__35127\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35568\,
            in1 => \N__42246\,
            in2 => \_gnd_net_\,
            in3 => \N__35106\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42038\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45141\,
            in1 => \N__42247\,
            in2 => \_gnd_net_\,
            in3 => \N__45105\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__42250\,
            in1 => \N__35274\,
            in2 => \N__35244\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45224\,
            in1 => \N__42251\,
            in2 => \_gnd_net_\,
            in3 => \N__45183\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46968\,
            in1 => \N__47350\,
            in2 => \N__44776\,
            in3 => \N__44733\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36750\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__42252\,
            in1 => \N__35193\,
            in2 => \N__35472\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__47351\,
            in1 => \N__46969\,
            in2 => \N__44952\,
            in3 => \N__44986\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42253\,
            in1 => \N__47439\,
            in2 => \_gnd_net_\,
            in3 => \N__47466\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44679\,
            in1 => \N__42254\,
            in2 => \_gnd_net_\,
            in3 => \N__44697\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37558\,
            in2 => \N__37495\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__46022\,
            ce => \N__41019\,
            sr => \N__45589\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38113\,
            in2 => \N__37528\,
            in3 => \N__35402\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__46022\,
            ce => \N__41019\,
            sr => \N__45589\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38089\,
            in2 => \N__37496\,
            in3 => \N__35351\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__46022\,
            ce => \N__41019\,
            sr => \N__45589\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38065\,
            in2 => \N__38117\,
            in3 => \N__35306\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__46022\,
            ce => \N__41019\,
            sr => \N__45589\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38090\,
            in2 => \N__38041\,
            in3 => \N__35303\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__46022\,
            ce => \N__41019\,
            sr => \N__45589\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38014\,
            in2 => \N__38069\,
            in3 => \N__35300\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__46022\,
            ce => \N__41019\,
            sr => \N__45589\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37990\,
            in2 => \N__38042\,
            in3 => \N__35297\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__46022\,
            ce => \N__41019\,
            sr => \N__45589\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38015\,
            in2 => \N__37966\,
            in3 => \N__35255\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__46022\,
            ce => \N__41019\,
            sr => \N__45589\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37936\,
            in2 => \N__37994\,
            in3 => \N__35534\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__46017\,
            ce => \N__41018\,
            sr => \N__45593\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38347\,
            in2 => \N__37967\,
            in3 => \N__35531\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__46017\,
            ce => \N__41018\,
            sr => \N__45593\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37937\,
            in2 => \N__38324\,
            in3 => \N__35528\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__46017\,
            ce => \N__41018\,
            sr => \N__45593\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38293\,
            in2 => \N__38351\,
            in3 => \N__35525\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__46017\,
            ce => \N__41018\,
            sr => \N__45593\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38323\,
            in2 => \N__38269\,
            in3 => \N__35522\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__46017\,
            ce => \N__41018\,
            sr => \N__45593\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38242\,
            in2 => \N__38297\,
            in3 => \N__35483\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__46017\,
            ce => \N__41018\,
            sr => \N__45593\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38218\,
            in2 => \N__38270\,
            in3 => \N__35480\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__46017\,
            ce => \N__41018\,
            sr => \N__45593\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38243\,
            in2 => \N__38195\,
            in3 => \N__35477\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__46017\,
            ce => \N__41018\,
            sr => \N__45593\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38161\,
            in2 => \N__38222\,
            in3 => \N__35444\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__46014\,
            ce => \N__41017\,
            sr => \N__45600\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38137\,
            in2 => \N__38194\,
            in3 => \N__35600\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__46014\,
            ce => \N__41017\,
            sr => \N__45600\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38162\,
            in2 => \N__38558\,
            in3 => \N__35597\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__46014\,
            ce => \N__41017\,
            sr => \N__45600\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38527\,
            in2 => \N__38141\,
            in3 => \N__35594\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__46014\,
            ce => \N__41017\,
            sr => \N__45600\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38557\,
            in2 => \N__38503\,
            in3 => \N__35591\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__46014\,
            ce => \N__41017\,
            sr => \N__45600\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38476\,
            in2 => \N__38531\,
            in3 => \N__35588\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__46014\,
            ce => \N__41017\,
            sr => \N__45600\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38452\,
            in2 => \N__38504\,
            in3 => \N__35585\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__46014\,
            ce => \N__41017\,
            sr => \N__45600\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38477\,
            in2 => \N__38428\,
            in3 => \N__35582\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__46014\,
            ce => \N__41017\,
            sr => \N__45600\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38398\,
            in2 => \N__38456\,
            in3 => \N__35579\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__46011\,
            ce => \N__41016\,
            sr => \N__45607\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38374\,
            in2 => \N__38429\,
            in3 => \N__35576\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__46011\,
            ce => \N__41016\,
            sr => \N__45607\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38399\,
            in2 => \N__38933\,
            in3 => \N__35846\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__46011\,
            ce => \N__41016\,
            sr => \N__45607\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38783\,
            in2 => \N__38378\,
            in3 => \N__35843\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__46011\,
            ce => \N__41016\,
            sr => \N__45607\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35840\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__41182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41850\,
            in2 => \_gnd_net_\,
            in3 => \N__41888\,
            lcout => \phase_controller_inst2.start_timer_hc_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35819\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__35744\,
            in1 => \N__46286\,
            in2 => \_gnd_net_\,
            in3 => \N__46351\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46107\,
            ce => 'H',
            sr => \N__45514\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__35743\,
            in1 => \N__46285\,
            in2 => \_gnd_net_\,
            in3 => \N__46350\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_435_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35742\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39063\,
            in1 => \N__39012\,
            in2 => \N__42842\,
            in3 => \N__42785\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36252\,
            in1 => \N__36198\,
            in2 => \N__36317\,
            in3 => \N__36363\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__36199\,
            in1 => \N__38623\,
            in2 => \N__38675\,
            in3 => \N__36253\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__35930\,
            in1 => \N__36364\,
            in2 => \N__35933\,
            in3 => \N__38636\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35860\,
            in2 => \_gnd_net_\,
            in3 => \N__39382\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39011\,
            in1 => \N__36309\,
            in2 => \N__42790\,
            in3 => \N__39062\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35890\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46098\,
            ce => \N__38694\,
            sr => \N__45527\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__43102\,
            in1 => \N__38674\,
            in2 => \N__35923\,
            in3 => \N__42993\,
            lcout => \elapsed_time_ns_1_RNIAE2591_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36145\,
            in2 => \N__38726\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__46093\,
            ce => \N__38696\,
            sr => \N__45529\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36124\,
            in2 => \N__35894\,
            in3 => \N__35849\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__46093\,
            ce => \N__38696\,
            sr => \N__45529\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36146\,
            in2 => \N__36104\,
            in3 => \N__36128\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__46093\,
            ce => \N__38696\,
            sr => \N__45529\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36125\,
            in2 => \N__36077\,
            in3 => \N__36107\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__46093\,
            ce => \N__38696\,
            sr => \N__45529\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36103\,
            in2 => \N__36049\,
            in3 => \N__36080\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__46093\,
            ce => \N__38696\,
            sr => \N__45529\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36076\,
            in2 => \N__36022\,
            in3 => \N__36053\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__46093\,
            ce => \N__38696\,
            sr => \N__45529\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35989\,
            in2 => \N__36050\,
            in3 => \N__36026\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__46093\,
            ce => \N__38696\,
            sr => \N__45529\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35956\,
            in2 => \N__36023\,
            in3 => \N__35999\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__46093\,
            ce => \N__38696\,
            sr => \N__45529\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36457\,
            in2 => \N__35996\,
            in3 => \N__35966\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__46086\,
            ce => \N__38697\,
            sr => \N__45533\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36433\,
            in2 => \N__35963\,
            in3 => \N__35936\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__46086\,
            ce => \N__38697\,
            sr => \N__45533\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36458\,
            in2 => \N__36410\,
            in3 => \N__36440\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__46086\,
            ce => \N__38697\,
            sr => \N__45533\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36382\,
            in2 => \N__36437\,
            in3 => \N__36413\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__46086\,
            ce => \N__38697\,
            sr => \N__45533\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36409\,
            in2 => \N__36340\,
            in3 => \N__36386\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__46086\,
            ce => \N__38697\,
            sr => \N__45533\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36383\,
            in2 => \N__36283\,
            in3 => \N__36344\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__46086\,
            ce => \N__38697\,
            sr => \N__45533\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36226\,
            in2 => \N__36341\,
            in3 => \N__36287\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__46086\,
            ce => \N__38697\,
            sr => \N__45533\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36169\,
            in2 => \N__36284\,
            in3 => \N__36236\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__46086\,
            ce => \N__38697\,
            sr => \N__45533\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36712\,
            in2 => \N__36233\,
            in3 => \N__36179\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__46079\,
            ce => \N__38698\,
            sr => \N__45539\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36691\,
            in2 => \N__36176\,
            in3 => \N__36149\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__46079\,
            ce => \N__38698\,
            sr => \N__45539\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36713\,
            in2 => \N__36671\,
            in3 => \N__36695\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__46079\,
            ce => \N__38698\,
            sr => \N__45539\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36692\,
            in2 => \N__36644\,
            in3 => \N__36674\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__46079\,
            ce => \N__38698\,
            sr => \N__45539\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36670\,
            in2 => \N__36616\,
            in3 => \N__36647\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__46079\,
            ce => \N__38698\,
            sr => \N__45539\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36643\,
            in2 => \N__36589\,
            in3 => \N__36620\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__46079\,
            ce => \N__38698\,
            sr => \N__45539\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36556\,
            in2 => \N__36617\,
            in3 => \N__36593\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__46079\,
            ce => \N__38698\,
            sr => \N__45539\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36523\,
            in2 => \N__36590\,
            in3 => \N__36566\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__46079\,
            ce => \N__38698\,
            sr => \N__45539\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36499\,
            in2 => \N__36563\,
            in3 => \N__36533\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__46072\,
            ce => \N__38699\,
            sr => \N__45543\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36835\,
            in2 => \N__36530\,
            in3 => \N__36503\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__46072\,
            ce => \N__38699\,
            sr => \N__45543\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36500\,
            in2 => \N__36482\,
            in3 => \N__36461\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__46072\,
            ce => \N__38699\,
            sr => \N__45543\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36854\,
            in2 => \N__36839\,
            in3 => \N__36815\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__46072\,
            ce => \N__38699\,
            sr => \N__45543\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36812\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46072\,
            ce => \N__38699\,
            sr => \N__45543\
        );

    \phase_controller_inst2.T45_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__36802\,
            in1 => \N__41972\,
            in2 => \_gnd_net_\,
            in3 => \N__46168\,
            lcout => \T45_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46067\,
            ce => 'H',
            sr => \N__45548\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__37762\,
            in1 => \N__36788\,
            in2 => \_gnd_net_\,
            in3 => \N__37247\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__44078\,
            in1 => \_gnd_net_\,
            in2 => \N__36791\,
            in3 => \N__37763\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41057\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46060\,
            ce => \N__41024\,
            sr => \N__45551\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__44459\,
            in1 => \N__36782\,
            in2 => \_gnd_net_\,
            in3 => \N__40928\,
            lcout => \current_shift_inst.control_input_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.N_1572_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47256\,
            in1 => \N__36772\,
            in2 => \N__46800\,
            in3 => \N__36734\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__40931\,
            in1 => \N__44630\,
            in2 => \_gnd_net_\,
            in3 => \N__37016\,
            lcout => \current_shift_inst.control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__37007\,
            in1 => \N__44399\,
            in2 => \_gnd_net_\,
            in3 => \N__40930\,
            lcout => \current_shift_inst.control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37033\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47257\,
            in1 => \N__42394\,
            in2 => \N__46801\,
            in3 => \N__36985\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__40932\,
            in1 => \N__44615\,
            in2 => \_gnd_net_\,
            in3 => \N__36950\,
            lcout => \current_shift_inst.control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_0_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36941\,
            in2 => \N__36934\,
            in3 => \N__36935\,
            lcout => \current_shift_inst.control_inputZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \current_shift_inst.control_input_1_cry_0\,
            clk => \N__46046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37292\,
            in3 => \N__36881\,
            lcout => \current_shift_inst.control_inputZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_0\,
            carryout => \current_shift_inst.control_input_1_cry_1\,
            clk => \N__46046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_2_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37253\,
            in2 => \_gnd_net_\,
            in3 => \N__36863\,
            lcout => \current_shift_inst.control_inputZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_1\,
            carryout => \current_shift_inst.control_input_1_cry_2\,
            clk => \N__46046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_3_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36860\,
            in2 => \_gnd_net_\,
            in3 => \N__37157\,
            lcout => \current_shift_inst.control_inputZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_2\,
            carryout => \current_shift_inst.control_input_1_cry_3\,
            clk => \N__46046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_4_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37154\,
            in2 => \_gnd_net_\,
            in3 => \N__37136\,
            lcout => \current_shift_inst.control_inputZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_3\,
            carryout => \current_shift_inst.control_input_1_cry_4\,
            clk => \N__46046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_5_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37133\,
            in2 => \_gnd_net_\,
            in3 => \N__37112\,
            lcout => \current_shift_inst.control_inputZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_4\,
            carryout => \current_shift_inst.control_input_1_cry_5\,
            clk => \N__46046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_6_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40979\,
            in2 => \_gnd_net_\,
            in3 => \N__37100\,
            lcout => \current_shift_inst.control_inputZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_5\,
            carryout => \current_shift_inst.control_input_1_cry_6\,
            clk => \N__46046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_7_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37277\,
            in2 => \_gnd_net_\,
            in3 => \N__37082\,
            lcout => \current_shift_inst.control_inputZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_6\,
            carryout => \current_shift_inst.control_input_1_cry_7\,
            clk => \N__46046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_8_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40958\,
            in2 => \_gnd_net_\,
            in3 => \N__37067\,
            lcout => \current_shift_inst.control_inputZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \current_shift_inst.control_input_1_cry_8\,
            clk => \N__46040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_9_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40877\,
            in2 => \_gnd_net_\,
            in3 => \N__37064\,
            lcout => \current_shift_inst.control_inputZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_8\,
            carryout => \current_shift_inst.control_input_1_cry_9\,
            clk => \N__46040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_10_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37265\,
            in2 => \_gnd_net_\,
            in3 => \N__37049\,
            lcout => \current_shift_inst.control_inputZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_9\,
            carryout => \current_shift_inst.control_input_1_cry_10\,
            clk => \N__46040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_11_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37046\,
            in2 => \_gnd_net_\,
            in3 => \N__37040\,
            lcout => \current_shift_inst.control_inputZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__37298\,
            in1 => \N__44438\,
            in2 => \_gnd_net_\,
            in3 => \N__40933\,
            lcout => \current_shift_inst.control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__40935\,
            in1 => \N__37283\,
            in2 => \_gnd_net_\,
            in3 => \N__44582\,
            lcout => \current_shift_inst.control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__37271\,
            in1 => \N__44516\,
            in2 => \_gnd_net_\,
            in3 => \N__40936\,
            lcout => \current_shift_inst.control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__40934\,
            in1 => \N__44411\,
            in2 => \_gnd_net_\,
            in3 => \N__37259\,
            lcout => \current_shift_inst.control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37240\,
            in2 => \N__37223\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37817\,
            in2 => \N__37202\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37190\,
            in2 => \N__37880\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37821\,
            in2 => \N__37178\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37373\,
            in2 => \N__37881\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37825\,
            in2 => \N__37361\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37346\,
            in2 => \N__37882\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37829\,
            in2 => \N__37334\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37842\,
            in2 => \N__42056\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37319\,
            in2 => \N__37886\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37830\,
            in2 => \N__37313\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37304\,
            in2 => \N__37883\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37834\,
            in2 => \N__42410\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37604\,
            in2 => \N__37884\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37838\,
            in2 => \N__37421\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37412\,
            in2 => \N__37885\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37887\,
            in2 => \N__37406\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41276\,
            in2 => \N__37912\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37891\,
            in2 => \N__37397\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37388\,
            in2 => \N__37913\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37895\,
            in2 => \N__37382\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37897\,
            in2 => \N__41069\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37896\,
            in2 => \N__42266\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37898\,
            in2 => \N__41270\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37899\,
            in2 => \N__37595\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37583\,
            in2 => \N__37914\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37903\,
            in2 => \N__37466\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37448\,
            in2 => \N__37915\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37907\,
            in2 => \N__41150\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37433\,
            in2 => \N__37916\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37911\,
            in2 => \N__37622\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47369\,
            in2 => \_gnd_net_\,
            in3 => \N__37607\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42255\,
            in1 => \N__45060\,
            in2 => \_gnd_net_\,
            in3 => \N__45037\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42256\,
            in1 => \N__44841\,
            in2 => \_gnd_net_\,
            in3 => \N__44818\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47368\,
            in1 => \N__44979\,
            in2 => \_gnd_net_\,
            in3 => \N__44953\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42311\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38909\,
            in1 => \N__37554\,
            in2 => \_gnd_net_\,
            in3 => \N__37535\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__46018\,
            ce => \N__38750\,
            sr => \N__45594\
        );

    \current_shift_inst.timer_s1.counter_1_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38905\,
            in1 => \N__37518\,
            in2 => \_gnd_net_\,
            in3 => \N__37499\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__46018\,
            ce => \N__38750\,
            sr => \N__45594\
        );

    \current_shift_inst.timer_s1.counter_2_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38910\,
            in1 => \N__37483\,
            in2 => \_gnd_net_\,
            in3 => \N__37469\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__46018\,
            ce => \N__38750\,
            sr => \N__45594\
        );

    \current_shift_inst.timer_s1.counter_3_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38906\,
            in1 => \N__38112\,
            in2 => \_gnd_net_\,
            in3 => \N__38093\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__46018\,
            ce => \N__38750\,
            sr => \N__45594\
        );

    \current_shift_inst.timer_s1.counter_4_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38911\,
            in1 => \N__38088\,
            in2 => \_gnd_net_\,
            in3 => \N__38072\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__46018\,
            ce => \N__38750\,
            sr => \N__45594\
        );

    \current_shift_inst.timer_s1.counter_5_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38907\,
            in1 => \N__38064\,
            in2 => \_gnd_net_\,
            in3 => \N__38045\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__46018\,
            ce => \N__38750\,
            sr => \N__45594\
        );

    \current_shift_inst.timer_s1.counter_6_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38912\,
            in1 => \N__38034\,
            in2 => \_gnd_net_\,
            in3 => \N__38018\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__46018\,
            ce => \N__38750\,
            sr => \N__45594\
        );

    \current_shift_inst.timer_s1.counter_7_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38908\,
            in1 => \N__38013\,
            in2 => \_gnd_net_\,
            in3 => \N__37997\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__46018\,
            ce => \N__38750\,
            sr => \N__45594\
        );

    \current_shift_inst.timer_s1.counter_8_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38900\,
            in1 => \N__37989\,
            in2 => \_gnd_net_\,
            in3 => \N__37970\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__46015\,
            ce => \N__38767\,
            sr => \N__45601\
        );

    \current_shift_inst.timer_s1.counter_9_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38904\,
            in1 => \N__37959\,
            in2 => \_gnd_net_\,
            in3 => \N__37940\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__46015\,
            ce => \N__38767\,
            sr => \N__45601\
        );

    \current_shift_inst.timer_s1.counter_10_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38897\,
            in1 => \N__37935\,
            in2 => \_gnd_net_\,
            in3 => \N__37919\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__46015\,
            ce => \N__38767\,
            sr => \N__45601\
        );

    \current_shift_inst.timer_s1.counter_11_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38901\,
            in1 => \N__38346\,
            in2 => \_gnd_net_\,
            in3 => \N__38327\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__46015\,
            ce => \N__38767\,
            sr => \N__45601\
        );

    \current_shift_inst.timer_s1.counter_12_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38898\,
            in1 => \N__38319\,
            in2 => \_gnd_net_\,
            in3 => \N__38300\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__46015\,
            ce => \N__38767\,
            sr => \N__45601\
        );

    \current_shift_inst.timer_s1.counter_13_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38902\,
            in1 => \N__38292\,
            in2 => \_gnd_net_\,
            in3 => \N__38273\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__46015\,
            ce => \N__38767\,
            sr => \N__45601\
        );

    \current_shift_inst.timer_s1.counter_14_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38899\,
            in1 => \N__38262\,
            in2 => \_gnd_net_\,
            in3 => \N__38246\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__46015\,
            ce => \N__38767\,
            sr => \N__45601\
        );

    \current_shift_inst.timer_s1.counter_15_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38903\,
            in1 => \N__38241\,
            in2 => \_gnd_net_\,
            in3 => \N__38225\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__46015\,
            ce => \N__38767\,
            sr => \N__45601\
        );

    \current_shift_inst.timer_s1.counter_16_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38869\,
            in1 => \N__38217\,
            in2 => \_gnd_net_\,
            in3 => \N__38198\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_16_24_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__46012\,
            ce => \N__38768\,
            sr => \N__45608\
        );

    \current_shift_inst.timer_s1.counter_17_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38873\,
            in1 => \N__38184\,
            in2 => \_gnd_net_\,
            in3 => \N__38165\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__46012\,
            ce => \N__38768\,
            sr => \N__45608\
        );

    \current_shift_inst.timer_s1.counter_18_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38870\,
            in1 => \N__38160\,
            in2 => \_gnd_net_\,
            in3 => \N__38144\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__46012\,
            ce => \N__38768\,
            sr => \N__45608\
        );

    \current_shift_inst.timer_s1.counter_19_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38874\,
            in1 => \N__38136\,
            in2 => \_gnd_net_\,
            in3 => \N__38561\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__46012\,
            ce => \N__38768\,
            sr => \N__45608\
        );

    \current_shift_inst.timer_s1.counter_20_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38871\,
            in1 => \N__38553\,
            in2 => \_gnd_net_\,
            in3 => \N__38534\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__46012\,
            ce => \N__38768\,
            sr => \N__45608\
        );

    \current_shift_inst.timer_s1.counter_21_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38875\,
            in1 => \N__38526\,
            in2 => \_gnd_net_\,
            in3 => \N__38507\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__46012\,
            ce => \N__38768\,
            sr => \N__45608\
        );

    \current_shift_inst.timer_s1.counter_22_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38872\,
            in1 => \N__38496\,
            in2 => \_gnd_net_\,
            in3 => \N__38480\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__46012\,
            ce => \N__38768\,
            sr => \N__45608\
        );

    \current_shift_inst.timer_s1.counter_23_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38876\,
            in1 => \N__38475\,
            in2 => \_gnd_net_\,
            in3 => \N__38459\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__46012\,
            ce => \N__38768\,
            sr => \N__45608\
        );

    \current_shift_inst.timer_s1.counter_24_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38865\,
            in1 => \N__38451\,
            in2 => \_gnd_net_\,
            in3 => \N__38432\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_16_25_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__46006\,
            ce => \N__38766\,
            sr => \N__45622\
        );

    \current_shift_inst.timer_s1.counter_25_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38877\,
            in1 => \N__38421\,
            in2 => \_gnd_net_\,
            in3 => \N__38402\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__46006\,
            ce => \N__38766\,
            sr => \N__45622\
        );

    \current_shift_inst.timer_s1.counter_26_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38866\,
            in1 => \N__38397\,
            in2 => \_gnd_net_\,
            in3 => \N__38381\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__46006\,
            ce => \N__38766\,
            sr => \N__45622\
        );

    \current_shift_inst.timer_s1.counter_27_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38878\,
            in1 => \N__38373\,
            in2 => \_gnd_net_\,
            in3 => \N__38354\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__46006\,
            ce => \N__38766\,
            sr => \N__45622\
        );

    \current_shift_inst.timer_s1.counter_28_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38867\,
            in1 => \N__38929\,
            in2 => \_gnd_net_\,
            in3 => \N__38915\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__46006\,
            ce => \N__38766\,
            sr => \N__45622\
        );

    \current_shift_inst.timer_s1.counter_29_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__38782\,
            in1 => \N__38868\,
            in2 => \_gnd_net_\,
            in3 => \N__38786\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46006\,
            ce => \N__38766\,
            sr => \N__45622\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38725\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46108\,
            ce => \N__38695\,
            sr => \N__45515\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38670\,
            in1 => \N__38619\,
            in2 => \N__38653\,
            in3 => \N__38635\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__38590\,
            in1 => \N__43141\,
            in2 => \N__38624\,
            in3 => \N__39109\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38606\,
            in3 => \N__42695\,
            lcout => \elapsed_time_ns_1_RNIRHL2M1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__42670\,
            in1 => \N__42614\,
            in2 => \N__42647\,
            in3 => \N__42632\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_381\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__43427\,
            in1 => \N__43378\,
            in2 => \N__38564\,
            in3 => \N__42581\,
            lcout => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\,
            ltout => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__39398\,
            in1 => \N__39308\,
            in2 => \N__39152\,
            in3 => \N__42962\,
            lcout => \elapsed_time_ns_1_RNIRAIF91_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__45716\,
            in1 => \N__43377\,
            in2 => \_gnd_net_\,
            in3 => \N__42580\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__43428\,
            in1 => \N__45717\,
            in2 => \N__39149\,
            in3 => \N__39146\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38992\,
            in1 => \N__39317\,
            in2 => \N__39040\,
            in3 => \N__42810\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__39064\,
            in1 => \N__39033\,
            in2 => \N__42596\,
            in3 => \N__38991\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_348_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39316\,
            in2 => \N__39020\,
            in3 => \N__39013\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__43099\,
            in1 => \N__39331\,
            in2 => \N__39231\,
            in3 => \N__42957\,
            lcout => \elapsed_time_ns_1_RNIR9HF91_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__38993\,
            in1 => \N__43101\,
            in2 => \N__42983\,
            in3 => \N__38981\,
            lcout => \elapsed_time_ns_1_RNIFJ2591_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__43100\,
            in1 => \N__38939\,
            in2 => \N__39293\,
            in3 => \N__42958\,
            lcout => \elapsed_time_ns_1_RNITCIF91_0_23\,
            ltout => \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42529\,
            in1 => \N__43240\,
            in2 => \N__39401\,
            in3 => \N__39397\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43204\,
            in1 => \N__43463\,
            in2 => \N__39386\,
            in3 => \N__40091\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__43107\,
            in1 => \N__39383\,
            in2 => \N__39363\,
            in3 => \N__42951\,
            lcout => \elapsed_time_ns_1_RNIDH2591_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39274\,
            in1 => \N__43351\,
            in2 => \N__39332\,
            in3 => \N__40039\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39169\,
            in1 => \N__43453\,
            in2 => \N__43306\,
            in3 => \N__43189\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42544\,
            in1 => \N__39304\,
            in2 => \N__43267\,
            in3 => \N__39286\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__43103\,
            in1 => \N__39252\,
            in2 => \N__42975\,
            in3 => \N__39275\,
            lcout => \elapsed_time_ns_1_RNIQ8HF91_0_11\,
            ltout => \elapsed_time_ns_1_RNIQ8HF91_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__40017\,
            in1 => \N__43323\,
            in2 => \N__39239\,
            in3 => \N__39216\,
            lcout => \phase_controller_inst1.stoper_tr.N_244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__39170\,
            in1 => \N__42950\,
            in2 => \N__43145\,
            in3 => \N__39158\,
            lcout => \elapsed_time_ns_1_RNI3JIF91_0_29\,
            ltout => \elapsed_time_ns_1_RNI3JIF91_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__42853\,
            in1 => \_gnd_net_\,
            in2 => \N__40094\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__39998\,
            in1 => \N__39899\,
            in2 => \N__40085\,
            in3 => \N__39716\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46087\,
            ce => \N__39597\,
            sr => \N__45534\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__43137\,
            in1 => \N__40040\,
            in2 => \N__42992\,
            in3 => \N__40024\,
            lcout => \elapsed_time_ns_1_RNISAHF91_0_13\,
            ltout => \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__39997\,
            in1 => \N__39898\,
            in2 => \N__39941\,
            in3 => \N__39715\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46087\,
            ce => \N__39597\,
            sr => \N__45534\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__39926\,
            in1 => \N__39897\,
            in2 => \_gnd_net_\,
            in3 => \N__39714\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46087\,
            ce => \N__39597\,
            sr => \N__45534\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_1_c_inv_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44122\,
            in1 => \N__39467\,
            in2 => \N__39455\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_2_c_inv_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39443\,
            in2 => \N__39431\,
            in3 => \N__40490\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_3_c_inv_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39422\,
            in2 => \N__39410\,
            in3 => \N__40472\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_4_c_inv_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40265\,
            in2 => \N__40253\,
            in3 => \N__40454\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_5_c_inv_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40244\,
            in2 => \N__40232\,
            in3 => \N__40745\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_6_c_inv_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40727\,
            in1 => \N__40223\,
            in2 => \N__40211\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_7_c_inv_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40202\,
            in2 => \N__40190\,
            in3 => \N__40709\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_8_c_inv_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40181\,
            in2 => \N__40169\,
            in3 => \N__40691\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_9_c_inv_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40157\,
            in2 => \N__40145\,
            in3 => \N__40673\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_10_c_inv_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40136\,
            in2 => \N__40124\,
            in3 => \N__40655\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_11_c_inv_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40115\,
            in2 => \N__40103\,
            in3 => \N__40637\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_12_c_inv_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40436\,
            in2 => \N__40424\,
            in3 => \N__40619\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_13_c_inv_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40415\,
            in2 => \N__40403\,
            in3 => \N__40601\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_14_c_inv_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40868\,
            in1 => \N__40394\,
            in2 => \N__40382\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_15_c_inv_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40370\,
            in2 => \N__40358\,
            in3 => \N__40850\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_16_c_inv_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40349\,
            in2 => \N__40337\,
            in3 => \N__40829\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_17_c_inv_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40328\,
            in2 => \N__40316\,
            in3 => \N__40811\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_18_c_inv_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40307\,
            in2 => \N__40295\,
            in3 => \N__40793\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_inv_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40286\,
            in2 => \N__40274\,
            in3 => \N__40772\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40583\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43496\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44139\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNILGTP_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43565\,
            in2 => \_gnd_net_\,
            in3 => \N__43608\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a3_1_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40551\,
            in2 => \_gnd_net_\,
            in3 => \N__43664\,
            lcout => state_ns_i_a3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40496\,
            in2 => \N__44123\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44256\,
            in1 => \N__40489\,
            in2 => \_gnd_net_\,
            in3 => \N__40475\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__46061\,
            ce => 'H',
            sr => \N__45552\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__44271\,
            in1 => \N__40471\,
            in2 => \N__43592\,
            in3 => \N__40457\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__46061\,
            ce => 'H',
            sr => \N__45552\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44257\,
            in1 => \N__40453\,
            in2 => \_gnd_net_\,
            in3 => \N__40439\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__46061\,
            ce => 'H',
            sr => \N__45552\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44272\,
            in1 => \N__40744\,
            in2 => \_gnd_net_\,
            in3 => \N__40730\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__46061\,
            ce => 'H',
            sr => \N__45552\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44258\,
            in1 => \N__40726\,
            in2 => \_gnd_net_\,
            in3 => \N__40712\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__46061\,
            ce => 'H',
            sr => \N__45552\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44273\,
            in1 => \N__40708\,
            in2 => \_gnd_net_\,
            in3 => \N__40694\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__46061\,
            ce => 'H',
            sr => \N__45552\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44259\,
            in1 => \N__40690\,
            in2 => \_gnd_net_\,
            in3 => \N__40676\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__46061\,
            ce => 'H',
            sr => \N__45552\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44267\,
            in1 => \N__40672\,
            in2 => \_gnd_net_\,
            in3 => \N__40658\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__46053\,
            ce => 'H',
            sr => \N__45556\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44260\,
            in1 => \N__40654\,
            in2 => \_gnd_net_\,
            in3 => \N__40640\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__46053\,
            ce => 'H',
            sr => \N__45556\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44264\,
            in1 => \N__40636\,
            in2 => \_gnd_net_\,
            in3 => \N__40622\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__46053\,
            ce => 'H',
            sr => \N__45556\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44261\,
            in1 => \N__40618\,
            in2 => \_gnd_net_\,
            in3 => \N__40604\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__46053\,
            ce => 'H',
            sr => \N__45556\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44265\,
            in1 => \N__40600\,
            in2 => \_gnd_net_\,
            in3 => \N__40586\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__46053\,
            ce => 'H',
            sr => \N__45556\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44262\,
            in1 => \N__40867\,
            in2 => \_gnd_net_\,
            in3 => \N__40853\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__46053\,
            ce => 'H',
            sr => \N__45556\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44266\,
            in1 => \N__40846\,
            in2 => \_gnd_net_\,
            in3 => \N__40832\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__46053\,
            ce => 'H',
            sr => \N__45556\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44263\,
            in1 => \N__40828\,
            in2 => \_gnd_net_\,
            in3 => \N__40814\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__46053\,
            ce => 'H',
            sr => \N__45556\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44268\,
            in1 => \N__40810\,
            in2 => \_gnd_net_\,
            in3 => \N__40796\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__46047\,
            ce => 'H',
            sr => \N__45560\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44270\,
            in1 => \N__40792\,
            in2 => \_gnd_net_\,
            in3 => \N__40778\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__46047\,
            ce => 'H',
            sr => \N__45560\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44269\,
            in1 => \N__40771\,
            in2 => \_gnd_net_\,
            in3 => \N__40775\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46047\,
            ce => 'H',
            sr => \N__45560\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47344\,
            in1 => \N__41197\,
            in2 => \N__46980\,
            in3 => \N__41167\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__41198\,
            in1 => \N__47345\,
            in2 => \N__41171\,
            in3 => \N__46922\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47341\,
            in1 => \N__41196\,
            in2 => \_gnd_net_\,
            in3 => \N__41166\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_1_11_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47346\,
            in2 => \_gnd_net_\,
            in3 => \N__46918\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47342\,
            in1 => \N__41116\,
            in2 => \N__46981\,
            in3 => \N__41086\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__41117\,
            in1 => \N__47343\,
            in2 => \N__41090\,
            in3 => \N__46926\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42190\,
            in1 => \N__41115\,
            in2 => \_gnd_net_\,
            in3 => \N__41085\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41052\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46041\,
            ce => \N__41023\,
            sr => \N__45564\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__44591\,
            in1 => \N__40991\,
            in2 => \_gnd_net_\,
            in3 => \N__40925\,
            lcout => \current_shift_inst.control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__40926\,
            in1 => \N__44558\,
            in2 => \_gnd_net_\,
            in3 => \N__40970\,
            lcout => \current_shift_inst.control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__40949\,
            in1 => \N__44549\,
            in2 => \_gnd_net_\,
            in3 => \N__40927\,
            lcout => \current_shift_inst.control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__47339\,
            in1 => \N__41786\,
            in2 => \N__41750\,
            in3 => \N__46972\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__41717\,
            in1 => \N__41609\,
            in2 => \N__41579\,
            in3 => \N__41373\,
            lcout => \elapsed_time_ns_1_RNI81DJ11_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__47338\,
            in1 => \N__46971\,
            in2 => \N__42446\,
            in3 => \N__42488\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46970\,
            in1 => \N__47340\,
            in2 => \N__41354\,
            in3 => \N__41303\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46984\,
            in1 => \N__47354\,
            in2 => \N__42122\,
            in3 => \N__42083\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42218\,
            in1 => \N__41226\,
            in2 => \_gnd_net_\,
            in3 => \N__41253\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44775\,
            in1 => \N__42219\,
            in2 => \_gnd_net_\,
            in3 => \N__44734\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__47355\,
            in1 => \N__46983\,
            in2 => \N__41260\,
            in3 => \N__41227\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46982\,
            in1 => \N__47356\,
            in2 => \N__42340\,
            in3 => \N__42291\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42217\,
            in1 => \N__42486\,
            in2 => \_gnd_net_\,
            in3 => \N__42441\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__42386\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42220\,
            in1 => \N__42330\,
            in2 => \_gnd_net_\,
            in3 => \N__42293\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__42216\,
            in1 => \N__42111\,
            in2 => \_gnd_net_\,
            in3 => \N__42082\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47353\,
            in1 => \N__42043\,
            in2 => \N__47005\,
            in3 => \N__42014\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.T01_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__41899\,
            in1 => \N__41986\,
            in2 => \_gnd_net_\,
            in3 => \N__41857\,
            lcout => \T01_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46026\,
            ce => 'H',
            sr => \N__45583\
        );

    \phase_controller_inst2.state_1_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__43748\,
            in1 => \N__41887\,
            in2 => \N__46221\,
            in3 => \N__41846\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46019\,
            ce => 'H',
            sr => \N__45595\
        );

    \phase_controller_inst2.T12_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__41797\,
            in1 => \N__46229\,
            in2 => \_gnd_net_\,
            in3 => \N__41858\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46013\,
            ce => 'H',
            sr => \N__45609\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__42838\,
            in1 => \N__42823\,
            in2 => \N__42794\,
            in3 => \N__42755\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__43426\,
            in1 => \N__42631\,
            in2 => \N__42749\,
            in3 => \N__42643\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__45714\,
            in1 => \N__42674\,
            in2 => \N__42659\,
            in3 => \N__42613\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42517\,
            in1 => \N__43228\,
            in2 => \N__42571\,
            in3 => \N__42656\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__42630\,
            in1 => \N__42612\,
            in2 => \N__42599\,
            in3 => \N__42595\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_359_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__43475\,
            in1 => \N__42956\,
            in2 => \N__42572\,
            in3 => \N__43140\,
            lcout => \elapsed_time_ns_1_RNI0GIF91_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__42942\,
            in1 => \N__42551\,
            in2 => \N__42533\,
            in3 => \N__43073\,
            lcout => \elapsed_time_ns_1_RNIUDIF91_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__42518\,
            in1 => \N__42494\,
            in2 => \N__43121\,
            in3 => \N__42940\,
            lcout => \elapsed_time_ns_1_RNIVEIF91_0_25\,
            ltout => \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43438\,
            in1 => \N__43279\,
            in2 => \N__43478\,
            in3 => \N__43474\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__43069\,
            in1 => \N__43457\,
            in2 => \N__42991\,
            in3 => \N__43439\,
            lcout => \elapsed_time_ns_1_RNI2IIF91_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__43429\,
            in1 => \N__45715\,
            in2 => \N__43385\,
            in3 => \N__43361\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\,
            ltout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__43070\,
            in1 => \N__43355\,
            in2 => \N__43340\,
            in3 => \N__43329\,
            lcout => \elapsed_time_ns_1_RNIP7HF91_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__42941\,
            in1 => \N__43071\,
            in2 => \N__43286\,
            in3 => \N__43307\,
            lcout => \elapsed_time_ns_1_RNI1HIF91_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__43072\,
            in1 => \N__43268\,
            in2 => \N__43244\,
            in3 => \N__42943\,
            lcout => \elapsed_time_ns_1_RNISBIF91_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__43139\,
            in1 => \N__43229\,
            in2 => \N__42982\,
            in3 => \N__43205\,
            lcout => \elapsed_time_ns_1_RNIQ9IF91_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__43193\,
            in1 => \N__43138\,
            in2 => \N__42857\,
            in3 => \N__42952\,
            lcout => \elapsed_time_ns_1_RNIRBJF91_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__43825\,
            in1 => \N__43763\,
            in2 => \_gnd_net_\,
            in3 => \N__43933\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43934\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46094\,
            ce => 'H',
            sr => \N__45530\
        );

    \phase_controller_inst1.stoper_hc.running_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000101110"
        )
    port map (
            in0 => \N__43762\,
            in1 => \N__43877\,
            in2 => \N__43835\,
            in3 => \N__43793\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46088\,
            ce => 'H',
            sr => \N__45535\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46233\,
            in2 => \_gnd_net_\,
            in3 => \N__43741\,
            lcout => \phase_controller_inst2.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__43700\,
            in1 => \N__43694\,
            in2 => \N__43679\,
            in3 => \N__43524\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46073\,
            ce => 'H',
            sr => \N__45544\
        );

    \phase_controller_inst2.stoper_tr.running_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111001001110"
        )
    port map (
            in0 => \N__43498\,
            in1 => \N__43538\,
            in2 => \N__43572\,
            in3 => \N__43612\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46073\,
            ce => 'H',
            sr => \N__45544\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__43525\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46073\,
            ce => 'H',
            sr => \N__45544\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLH1_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43497\,
            in2 => \_gnd_net_\,
            in3 => \N__44140\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLHZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__43561\,
            in1 => \N__43537\,
            in2 => \_gnd_net_\,
            in3 => \N__43523\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__44243\,
            in1 => \N__44141\,
            in2 => \N__44126\,
            in3 => \N__44121\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46073\,
            ce => 'H',
            sr => \N__45544\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44099\,
            in2 => \N__44077\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44044\,
            in2 => \N__44021\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46651\,
            in2 => \N__44003\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43988\,
            in2 => \N__46824\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46655\,
            in2 => \N__43976\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43961\,
            in2 => \N__46825\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46659\,
            in2 => \N__43946\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44384\,
            in2 => \N__46826\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46827\,
            in2 => \N__44375\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44360\,
            in2 => \N__46957\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46831\,
            in2 => \N__44348\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45089\,
            in2 => \N__46958\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46835\,
            in2 => \N__44336\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45005\,
            in2 => \N__46959\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46839\,
            in2 => \N__44321\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44306\,
            in2 => \N__46960\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46843\,
            in2 => \N__45167\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44486\,
            in2 => \N__46961\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46847\,
            in2 => \N__44477\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47411\,
            in2 => \N__46962\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46851\,
            in2 => \N__44645\,
            in3 => \N__44447\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44444\,
            in2 => \N__46963\,
            in3 => \N__44429\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46855\,
            in2 => \N__44426\,
            in3 => \N__44402\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44714\,
            in2 => \N__46964\,
            in3 => \N__44387\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46859\,
            in2 => \N__44792\,
            in3 => \N__44618\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44927\,
            in2 => \N__46965\,
            in3 => \N__44603\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46863\,
            in2 => \N__44600\,
            in3 => \N__44585\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46364\,
            in2 => \N__46966\,
            in3 => \N__44570\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46867\,
            in2 => \N__44567\,
            in3 => \N__44552\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44864\,
            in2 => \N__46967\,
            in3 => \N__44543\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46871\,
            in2 => \N__44540\,
            in3 => \N__44504\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_2_11_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__46872\,
            in1 => \N__47367\,
            in2 => \_gnd_net_\,
            in3 => \N__44501\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46877\,
            in1 => \N__47364\,
            in2 => \N__45238\,
            in3 => \N__45191\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__47362\,
            in1 => \N__46875\,
            in2 => \N__45155\,
            in3 => \N__45113\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__46876\,
            in1 => \N__45079\,
            in2 => \N__45041\,
            in3 => \N__47363\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__47365\,
            in1 => \N__46874\,
            in2 => \N__44996\,
            in3 => \N__44957\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46873\,
            in1 => \N__47366\,
            in2 => \N__44921\,
            in3 => \N__44885\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46987\,
            in1 => \N__47360\,
            in2 => \N__44858\,
            in3 => \N__44819\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46985\,
            in1 => \N__47359\,
            in2 => \N__44780\,
            in3 => \N__44735\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__47358\,
            in1 => \N__46986\,
            in2 => \N__44705\,
            in3 => \N__44681\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__46988\,
            in1 => \N__47357\,
            in2 => \N__47474\,
            in3 => \N__47449\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47399\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47361\,
            in1 => \N__47047\,
            in2 => \N__47006\,
            in3 => \N__46393\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_18_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46273\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46256\,
            ce => 'H',
            sr => \N__45610\
        );

    \delay_measurement_inst.start_timer_tr_LC_18_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46272\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46256\,
            ce => 'H',
            sr => \N__45610\
        );

    \phase_controller_inst2.T23_LC_18_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__46129\,
            in1 => \N__46228\,
            in2 => \_gnd_net_\,
            in3 => \N__46175\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46007\,
            ce => 'H',
            sr => \N__45623\
        );
end \INTERFACE\;
