-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jul 10 2025 20:22:24

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__50761\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50759\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50748\ : std_logic;
signal \N__50741\ : std_logic;
signal \N__50740\ : std_logic;
signal \N__50739\ : std_logic;
signal \N__50732\ : std_logic;
signal \N__50731\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50723\ : std_logic;
signal \N__50722\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50714\ : std_logic;
signal \N__50713\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50705\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50703\ : std_logic;
signal \N__50696\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50687\ : std_logic;
signal \N__50686\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50677\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50668\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50658\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50650\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50632\ : std_logic;
signal \N__50631\ : std_logic;
signal \N__50628\ : std_logic;
signal \N__50625\ : std_logic;
signal \N__50624\ : std_logic;
signal \N__50619\ : std_logic;
signal \N__50616\ : std_logic;
signal \N__50613\ : std_logic;
signal \N__50608\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50598\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50592\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50577\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50570\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50550\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50531\ : std_logic;
signal \N__50530\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50522\ : std_logic;
signal \N__50521\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50519\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50511\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50504\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50383\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50249\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50246\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50235\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50232\ : std_logic;
signal \N__50231\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50229\ : std_logic;
signal \N__50228\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50225\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50222\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50216\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50213\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50211\ : std_logic;
signal \N__50210\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50207\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50204\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50196\ : std_logic;
signal \N__50195\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50193\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50190\ : std_logic;
signal \N__50189\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50186\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50167\ : std_logic;
signal \N__50166\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50163\ : std_logic;
signal \N__50162\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50159\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50156\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50149\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50146\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50139\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50136\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50133\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50130\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50127\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49814\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49788\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49728\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49725\ : std_logic;
signal \N__49724\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49722\ : std_logic;
signal \N__49721\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49694\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49689\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49676\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49673\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49670\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49668\ : std_logic;
signal \N__49667\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49664\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49662\ : std_logic;
signal \N__49661\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49654\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49647\ : std_logic;
signal \N__49646\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49644\ : std_logic;
signal \N__49643\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49641\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49637\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49632\ : std_logic;
signal \N__49631\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49622\ : std_logic;
signal \N__49621\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49613\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49607\ : std_logic;
signal \N__49604\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49284\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49278\ : std_logic;
signal \N__49275\ : std_logic;
signal \N__49274\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49258\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49251\ : std_logic;
signal \N__49248\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49228\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49206\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49174\ : std_logic;
signal \N__49171\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49139\ : std_logic;
signal \N__49134\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49085\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49062\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49052\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49002\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48996\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48960\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48951\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48918\ : std_logic;
signal \N__48915\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48906\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48824\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48810\ : std_logic;
signal \N__48807\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48726\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48630\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48612\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48560\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48515\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48499\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48485\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48374\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48356\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48271\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48058\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48019\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48005\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47952\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47338\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47251\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47219\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47108\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47035\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47023\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46774\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46753\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46705\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46636\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46283\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45918\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45898\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45817\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45703\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45351\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45068\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44380\ : std_logic;
signal \N__44377\ : std_logic;
signal \N__44374\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43782\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43738\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43535\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42457\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41680\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41398\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41392\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41048\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40042\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal \N_34_i_i\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_9 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \current_shift_inst.PI_CTRL.N_164\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_164_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_120\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_167\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_168\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_166\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \rgb_drv_RNOZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_162\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal \bfn_3_8_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.state_RNI7NN7Z0Z_0\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_302_i\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_\ : std_logic;
signal state_ns_i_a3_1 : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal s4_phy_c : std_logic;
signal il_max_comp1_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_53\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal s3_phy_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \delay_measurement_inst.hc_stateZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_26\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_248\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_248_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_55\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\ : std_logic;
signal \bfn_10_25_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\ : std_logic;
signal \bfn_10_26_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\ : std_logic;
signal delay_hc_input_c : std_logic;
signal delay_hc_d1 : std_logic;
signal delay_hc_d2 : std_logic;
signal \delay_measurement_inst.prev_hc_sigZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal measured_delay_tr_7 : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal measured_delay_tr_8 : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal measured_delay_tr_5 : std_logic;
signal measured_delay_tr_4 : std_logic;
signal measured_delay_tr_9 : std_logic;
signal measured_delay_tr_3 : std_logic;
signal measured_delay_tr_2 : std_logic;
signal measured_delay_tr_6 : std_logic;
signal measured_delay_tr_1 : std_logic;
signal measured_delay_tr_14 : std_logic;
signal measured_delay_tr_12 : std_logic;
signal measured_delay_tr_11 : std_logic;
signal measured_delay_tr_13 : std_logic;
signal measured_delay_tr_10 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\ : std_logic;
signal measured_delay_tr_16 : std_logic;
signal \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_RNO_0_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_72\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \delay_measurement_inst.N_267\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_287_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_290\ : std_logic;
signal \delay_measurement_inst.N_59\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_\ : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i\ : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7\ : std_logic;
signal \delay_measurement_inst.N_299\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_287_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\ : std_logic;
signal \delay_measurement_inst.N_265\ : std_logic;
signal \delay_measurement_inst.N_265_cascade_\ : std_logic;
signal \delay_measurement_inst.N_270\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\ : std_logic;
signal measured_delay_tr_17 : std_logic;
signal measured_delay_tr_18 : std_logic;
signal \delay_measurement_inst.N_325\ : std_logic;
signal measured_delay_tr_19 : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlt31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt9_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt31_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal measured_delay_hc_10 : std_logic;
signal measured_delay_hc_31 : std_logic;
signal measured_delay_hc_3 : std_logic;
signal measured_delay_hc_12 : std_logic;
signal measured_delay_hc_18 : std_logic;
signal measured_delay_hc_17 : std_logic;
signal measured_delay_hc_5 : std_logic;
signal measured_delay_hc_11 : std_logic;
signal measured_delay_hc_9 : std_logic;
signal measured_delay_hc_14 : std_logic;
signal measured_delay_hc_6 : std_logic;
signal measured_delay_hc_13 : std_logic;
signal measured_delay_hc_24 : std_logic;
signal measured_delay_hc_25 : std_logic;
signal measured_delay_hc_26 : std_logic;
signal measured_delay_hc_23 : std_logic;
signal state_3 : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_enablelt3_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_71\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_15\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_23\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_8\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_16\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlt3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\ : std_logic;
signal measured_delay_hc_22 : std_logic;
signal measured_delay_hc_7 : std_logic;
signal measured_delay_hc_0 : std_logic;
signal measured_delay_hc_20 : std_logic;
signal measured_delay_hc_16 : std_logic;
signal measured_delay_hc_1 : std_logic;
signal measured_delay_hc_8 : std_logic;
signal measured_delay_hc_21 : std_logic;
signal measured_delay_hc_15 : std_logic;
signal measured_delay_hc_4 : std_logic;
signal measured_delay_hc_2 : std_logic;
signal measured_delay_hc_19 : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt19_0_cascade_\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.N_180_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\ : std_logic;
signal measured_delay_tr_15 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_0\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_1_cry_0\ : std_logic;
signal \current_shift_inst.control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_8\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_13\ : std_logic;
signal \current_shift_inst.control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_14\ : std_logic;
signal \current_shift_inst.control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_15\ : std_logic;
signal \current_shift_inst.control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_16\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_17\ : std_logic;
signal \current_shift_inst.control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_18\ : std_logic;
signal \current_shift_inst.control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_19\ : std_logic;
signal \current_shift_inst.control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_20\ : std_logic;
signal \current_shift_inst.control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_21\ : std_logic;
signal \current_shift_inst.control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_22\ : std_logic;
signal \current_shift_inst.control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_23\ : std_logic;
signal \current_shift_inst.control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_24\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.N_1355_i\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_6\ : std_logic;
signal \current_shift_inst.control_input_1_axb_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_7\ : std_logic;
signal \current_shift_inst.control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \current_shift_inst.control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_303_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_3\ : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_11\ : std_logic;
signal \bfn_14_27_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_14_28_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_14_29_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal delay_tr_input_c : std_logic;
signal delay_tr_d1 : std_logic;
signal red_c_i : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_3\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_11\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_19\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_8\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_16\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_302_i_g\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_304_i\ : std_logic;
signal \delay_measurement_inst.tr_stateZ0Z_0\ : std_logic;
signal delay_tr_d2 : std_logic;
signal \delay_measurement_inst.prev_tr_sigZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_26\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI4Q3UZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI8V4UZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIC46UZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIG97UZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIKE8UZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIOJ9UZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIA1B41Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIL0S01Z0Z_11\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIP5T01Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNITAU01Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNICE9PZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIGJAPZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIS2EPZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIENGPZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIDGBQZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIHLCQZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8JZ0\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5KZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_30\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_0_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNICIEQZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.un4_control_input_0_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_17\ : std_logic;
signal measured_delay_hc_29 : std_logic;
signal measured_delay_hc_30 : std_logic;
signal measured_delay_hc_27 : std_logic;
signal \delay_measurement_inst.un1_elapsed_time_hc\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3\ : std_logic;
signal measured_delay_hc_28 : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIOTCPZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIGNFQZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI9BAQZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_12\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_305_i\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIKOBPZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI898PZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_11\ : std_logic;
signal \current_shift_inst.control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_13\ : std_logic;
signal \current_shift_inst.control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_18_21_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_180_i_g\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_18_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_18_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_18_24_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_18_25_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_181_i_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_304_i_g\ : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21505\&\N__21508\&\N__21506\&\N__21509\&\N__21507\&\N__19943\&\N__19966\&\N__20000\&\N__19925\&\N__19987\&\N__20902\&\N__20933\&\N__20020\&\N__20035\&\N__20050\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__38394\&\N__38391\&'0'&'0'&'0'&\N__38389\&\N__38393\&\N__38390\&\N__38392\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21608\&\N__21600\&\N__21606\&\N__21599\&\N__21607\&\N__21598\&\N__21609\&\N__21595\&\N__21602\&\N__21594\&\N__21603\&\N__21596\&\N__21604\&\N__21597\&\N__21605\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__38368\&\N__38365\&'0'&'0'&'0'&\N__38363\&\N__38367\&\N__38364\&\N__38366\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__23836\,
            RESETB => \N__36395\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__38398\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__38388\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__38279\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__38362\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__50759\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50761\,
            DIN => \N__50760\,
            DOUT => \N__50759\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50761\,
            PADOUT => \N__50760\,
            PADIN => \N__50759\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50750\,
            DIN => \N__50749\,
            DOUT => \N__50748\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50750\,
            PADOUT => \N__50749\,
            PADIN => \N__50748\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22012\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50741\,
            DIN => \N__50740\,
            DOUT => \N__50739\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50741\,
            PADOUT => \N__50740\,
            PADIN => \N__50739\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50732\,
            DIN => \N__50731\,
            DOUT => \N__50730\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50732\,
            PADOUT => \N__50731\,
            PADIN => \N__50730\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26020\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50723\,
            DIN => \N__50722\,
            DOUT => \N__50721\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50723\,
            PADOUT => \N__50722\,
            PADIN => \N__50721\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50714\,
            DIN => \N__50713\,
            DOUT => \N__50712\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50714\,
            PADOUT => \N__50713\,
            PADIN => \N__50712\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50705\,
            DIN => \N__50704\,
            DOUT => \N__50703\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50705\,
            PADOUT => \N__50704\,
            PADIN => \N__50703\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50696\,
            DIN => \N__50695\,
            DOUT => \N__50694\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50696\,
            PADOUT => \N__50695\,
            PADIN => \N__50694\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32089\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50687\,
            DIN => \N__50686\,
            DOUT => \N__50685\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50687\,
            PADOUT => \N__50686\,
            PADIN => \N__50685\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50678\,
            DIN => \N__50677\,
            DOUT => \N__50676\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50678\,
            PADOUT => \N__50677\,
            PADIN => \N__50676\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50669\,
            DIN => \N__50668\,
            DOUT => \N__50667\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50669\,
            PADOUT => \N__50668\,
            PADIN => \N__50667\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26071\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50660\,
            DIN => \N__50659\,
            DOUT => \N__50658\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50660\,
            PADOUT => \N__50659\,
            PADIN => \N__50658\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50651\,
            DIN => \N__50650\,
            DOUT => \N__50649\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50651\,
            PADOUT => \N__50650\,
            PADIN => \N__50649\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11973\ : InMux
    port map (
            O => \N__50632\,
            I => \N__50628\
        );

    \I__11972\ : InMux
    port map (
            O => \N__50631\,
            I => \N__50625\
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__50628\,
            I => \N__50619\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__50625\,
            I => \N__50619\
        );

    \I__11969\ : InMux
    port map (
            O => \N__50624\,
            I => \N__50616\
        );

    \I__11968\ : Span4Mux_v
    port map (
            O => \N__50619\,
            I => \N__50613\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__50616\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__11966\ : Odrv4
    port map (
            O => \N__50613\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__11965\ : InMux
    port map (
            O => \N__50608\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__11964\ : CascadeMux
    port map (
            O => \N__50605\,
            I => \N__50601\
        );

    \I__11963\ : CascadeMux
    port map (
            O => \N__50604\,
            I => \N__50598\
        );

    \I__11962\ : InMux
    port map (
            O => \N__50601\,
            I => \N__50592\
        );

    \I__11961\ : InMux
    port map (
            O => \N__50598\,
            I => \N__50592\
        );

    \I__11960\ : InMux
    port map (
            O => \N__50597\,
            I => \N__50589\
        );

    \I__11959\ : LocalMux
    port map (
            O => \N__50592\,
            I => \N__50586\
        );

    \I__11958\ : LocalMux
    port map (
            O => \N__50589\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__11957\ : Odrv12
    port map (
            O => \N__50586\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__11956\ : InMux
    port map (
            O => \N__50581\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__11955\ : CascadeMux
    port map (
            O => \N__50578\,
            I => \N__50574\
        );

    \I__11954\ : CascadeMux
    port map (
            O => \N__50577\,
            I => \N__50571\
        );

    \I__11953\ : InMux
    port map (
            O => \N__50574\,
            I => \N__50565\
        );

    \I__11952\ : InMux
    port map (
            O => \N__50571\,
            I => \N__50565\
        );

    \I__11951\ : InMux
    port map (
            O => \N__50570\,
            I => \N__50562\
        );

    \I__11950\ : LocalMux
    port map (
            O => \N__50565\,
            I => \N__50559\
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__50562\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__11948\ : Odrv12
    port map (
            O => \N__50559\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__11947\ : InMux
    port map (
            O => \N__50554\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__11946\ : InMux
    port map (
            O => \N__50551\,
            I => \N__50547\
        );

    \I__11945\ : InMux
    port map (
            O => \N__50550\,
            I => \N__50544\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__50547\,
            I => \N__50541\
        );

    \I__11943\ : LocalMux
    port map (
            O => \N__50544\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__11942\ : Odrv12
    port map (
            O => \N__50541\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__11941\ : InMux
    port map (
            O => \N__50536\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__11940\ : InMux
    port map (
            O => \N__50533\,
            I => \N__50499\
        );

    \I__11939\ : InMux
    port map (
            O => \N__50532\,
            I => \N__50499\
        );

    \I__11938\ : InMux
    port map (
            O => \N__50531\,
            I => \N__50490\
        );

    \I__11937\ : InMux
    port map (
            O => \N__50530\,
            I => \N__50490\
        );

    \I__11936\ : InMux
    port map (
            O => \N__50529\,
            I => \N__50490\
        );

    \I__11935\ : InMux
    port map (
            O => \N__50528\,
            I => \N__50490\
        );

    \I__11934\ : InMux
    port map (
            O => \N__50527\,
            I => \N__50481\
        );

    \I__11933\ : InMux
    port map (
            O => \N__50526\,
            I => \N__50481\
        );

    \I__11932\ : InMux
    port map (
            O => \N__50525\,
            I => \N__50481\
        );

    \I__11931\ : InMux
    port map (
            O => \N__50524\,
            I => \N__50481\
        );

    \I__11930\ : InMux
    port map (
            O => \N__50523\,
            I => \N__50472\
        );

    \I__11929\ : InMux
    port map (
            O => \N__50522\,
            I => \N__50472\
        );

    \I__11928\ : InMux
    port map (
            O => \N__50521\,
            I => \N__50472\
        );

    \I__11927\ : InMux
    port map (
            O => \N__50520\,
            I => \N__50472\
        );

    \I__11926\ : InMux
    port map (
            O => \N__50519\,
            I => \N__50463\
        );

    \I__11925\ : InMux
    port map (
            O => \N__50518\,
            I => \N__50463\
        );

    \I__11924\ : InMux
    port map (
            O => \N__50517\,
            I => \N__50463\
        );

    \I__11923\ : InMux
    port map (
            O => \N__50516\,
            I => \N__50463\
        );

    \I__11922\ : InMux
    port map (
            O => \N__50515\,
            I => \N__50454\
        );

    \I__11921\ : InMux
    port map (
            O => \N__50514\,
            I => \N__50454\
        );

    \I__11920\ : InMux
    port map (
            O => \N__50513\,
            I => \N__50454\
        );

    \I__11919\ : InMux
    port map (
            O => \N__50512\,
            I => \N__50454\
        );

    \I__11918\ : InMux
    port map (
            O => \N__50511\,
            I => \N__50445\
        );

    \I__11917\ : InMux
    port map (
            O => \N__50510\,
            I => \N__50445\
        );

    \I__11916\ : InMux
    port map (
            O => \N__50509\,
            I => \N__50445\
        );

    \I__11915\ : InMux
    port map (
            O => \N__50508\,
            I => \N__50445\
        );

    \I__11914\ : InMux
    port map (
            O => \N__50507\,
            I => \N__50436\
        );

    \I__11913\ : InMux
    port map (
            O => \N__50506\,
            I => \N__50436\
        );

    \I__11912\ : InMux
    port map (
            O => \N__50505\,
            I => \N__50436\
        );

    \I__11911\ : InMux
    port map (
            O => \N__50504\,
            I => \N__50436\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__50499\,
            I => \N__50427\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__50490\,
            I => \N__50427\
        );

    \I__11908\ : LocalMux
    port map (
            O => \N__50481\,
            I => \N__50427\
        );

    \I__11907\ : LocalMux
    port map (
            O => \N__50472\,
            I => \N__50427\
        );

    \I__11906\ : LocalMux
    port map (
            O => \N__50463\,
            I => \N__50418\
        );

    \I__11905\ : LocalMux
    port map (
            O => \N__50454\,
            I => \N__50418\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__50445\,
            I => \N__50418\
        );

    \I__11903\ : LocalMux
    port map (
            O => \N__50436\,
            I => \N__50418\
        );

    \I__11902\ : Span4Mux_v
    port map (
            O => \N__50427\,
            I => \N__50413\
        );

    \I__11901\ : Span4Mux_v
    port map (
            O => \N__50418\,
            I => \N__50413\
        );

    \I__11900\ : Odrv4
    port map (
            O => \N__50413\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__11899\ : InMux
    port map (
            O => \N__50410\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__11898\ : InMux
    port map (
            O => \N__50407\,
            I => \N__50404\
        );

    \I__11897\ : LocalMux
    port map (
            O => \N__50404\,
            I => \N__50400\
        );

    \I__11896\ : InMux
    port map (
            O => \N__50403\,
            I => \N__50397\
        );

    \I__11895\ : Span4Mux_h
    port map (
            O => \N__50400\,
            I => \N__50394\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__50397\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__11893\ : Odrv4
    port map (
            O => \N__50394\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__11892\ : CEMux
    port map (
            O => \N__50389\,
            I => \N__50386\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__50386\,
            I => \N__50380\
        );

    \I__11890\ : CEMux
    port map (
            O => \N__50385\,
            I => \N__50377\
        );

    \I__11889\ : CEMux
    port map (
            O => \N__50384\,
            I => \N__50374\
        );

    \I__11888\ : CEMux
    port map (
            O => \N__50383\,
            I => \N__50371\
        );

    \I__11887\ : Span4Mux_v
    port map (
            O => \N__50380\,
            I => \N__50368\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__50377\,
            I => \N__50365\
        );

    \I__11885\ : LocalMux
    port map (
            O => \N__50374\,
            I => \N__50362\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__50371\,
            I => \N__50359\
        );

    \I__11883\ : Span4Mux_h
    port map (
            O => \N__50368\,
            I => \N__50354\
        );

    \I__11882\ : Span4Mux_v
    port map (
            O => \N__50365\,
            I => \N__50354\
        );

    \I__11881\ : Span4Mux_h
    port map (
            O => \N__50362\,
            I => \N__50351\
        );

    \I__11880\ : Span4Mux_h
    port map (
            O => \N__50359\,
            I => \N__50348\
        );

    \I__11879\ : Span4Mux_h
    port map (
            O => \N__50354\,
            I => \N__50345\
        );

    \I__11878\ : Span4Mux_h
    port map (
            O => \N__50351\,
            I => \N__50342\
        );

    \I__11877\ : Span4Mux_h
    port map (
            O => \N__50348\,
            I => \N__50339\
        );

    \I__11876\ : Odrv4
    port map (
            O => \N__50345\,
            I => \current_shift_inst.timer_s1.N_181_i_g\
        );

    \I__11875\ : Odrv4
    port map (
            O => \N__50342\,
            I => \current_shift_inst.timer_s1.N_181_i_g\
        );

    \I__11874\ : Odrv4
    port map (
            O => \N__50339\,
            I => \current_shift_inst.timer_s1.N_181_i_g\
        );

    \I__11873\ : InMux
    port map (
            O => \N__50332\,
            I => \N__50329\
        );

    \I__11872\ : LocalMux
    port map (
            O => \N__50329\,
            I => \N__50325\
        );

    \I__11871\ : InMux
    port map (
            O => \N__50328\,
            I => \N__50322\
        );

    \I__11870\ : Span4Mux_h
    port map (
            O => \N__50325\,
            I => \N__50318\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__50322\,
            I => \N__50315\
        );

    \I__11868\ : InMux
    port map (
            O => \N__50321\,
            I => \N__50312\
        );

    \I__11867\ : Odrv4
    port map (
            O => \N__50318\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__11866\ : Odrv4
    port map (
            O => \N__50315\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__11865\ : LocalMux
    port map (
            O => \N__50312\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__11864\ : InMux
    port map (
            O => \N__50305\,
            I => \N__50301\
        );

    \I__11863\ : CascadeMux
    port map (
            O => \N__50304\,
            I => \N__50298\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__50301\,
            I => \N__50295\
        );

    \I__11861\ : InMux
    port map (
            O => \N__50298\,
            I => \N__50292\
        );

    \I__11860\ : Span4Mux_v
    port map (
            O => \N__50295\,
            I => \N__50287\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__50292\,
            I => \N__50287\
        );

    \I__11858\ : Span4Mux_h
    port map (
            O => \N__50287\,
            I => \N__50284\
        );

    \I__11857\ : Span4Mux_h
    port map (
            O => \N__50284\,
            I => \N__50281\
        );

    \I__11856\ : Odrv4
    port map (
            O => \N__50281\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__11855\ : ClkMux
    port map (
            O => \N__50278\,
            I => \N__49819\
        );

    \I__11854\ : ClkMux
    port map (
            O => \N__50277\,
            I => \N__49819\
        );

    \I__11853\ : ClkMux
    port map (
            O => \N__50276\,
            I => \N__49819\
        );

    \I__11852\ : ClkMux
    port map (
            O => \N__50275\,
            I => \N__49819\
        );

    \I__11851\ : ClkMux
    port map (
            O => \N__50274\,
            I => \N__49819\
        );

    \I__11850\ : ClkMux
    port map (
            O => \N__50273\,
            I => \N__49819\
        );

    \I__11849\ : ClkMux
    port map (
            O => \N__50272\,
            I => \N__49819\
        );

    \I__11848\ : ClkMux
    port map (
            O => \N__50271\,
            I => \N__49819\
        );

    \I__11847\ : ClkMux
    port map (
            O => \N__50270\,
            I => \N__49819\
        );

    \I__11846\ : ClkMux
    port map (
            O => \N__50269\,
            I => \N__49819\
        );

    \I__11845\ : ClkMux
    port map (
            O => \N__50268\,
            I => \N__49819\
        );

    \I__11844\ : ClkMux
    port map (
            O => \N__50267\,
            I => \N__49819\
        );

    \I__11843\ : ClkMux
    port map (
            O => \N__50266\,
            I => \N__49819\
        );

    \I__11842\ : ClkMux
    port map (
            O => \N__50265\,
            I => \N__49819\
        );

    \I__11841\ : ClkMux
    port map (
            O => \N__50264\,
            I => \N__49819\
        );

    \I__11840\ : ClkMux
    port map (
            O => \N__50263\,
            I => \N__49819\
        );

    \I__11839\ : ClkMux
    port map (
            O => \N__50262\,
            I => \N__49819\
        );

    \I__11838\ : ClkMux
    port map (
            O => \N__50261\,
            I => \N__49819\
        );

    \I__11837\ : ClkMux
    port map (
            O => \N__50260\,
            I => \N__49819\
        );

    \I__11836\ : ClkMux
    port map (
            O => \N__50259\,
            I => \N__49819\
        );

    \I__11835\ : ClkMux
    port map (
            O => \N__50258\,
            I => \N__49819\
        );

    \I__11834\ : ClkMux
    port map (
            O => \N__50257\,
            I => \N__49819\
        );

    \I__11833\ : ClkMux
    port map (
            O => \N__50256\,
            I => \N__49819\
        );

    \I__11832\ : ClkMux
    port map (
            O => \N__50255\,
            I => \N__49819\
        );

    \I__11831\ : ClkMux
    port map (
            O => \N__50254\,
            I => \N__49819\
        );

    \I__11830\ : ClkMux
    port map (
            O => \N__50253\,
            I => \N__49819\
        );

    \I__11829\ : ClkMux
    port map (
            O => \N__50252\,
            I => \N__49819\
        );

    \I__11828\ : ClkMux
    port map (
            O => \N__50251\,
            I => \N__49819\
        );

    \I__11827\ : ClkMux
    port map (
            O => \N__50250\,
            I => \N__49819\
        );

    \I__11826\ : ClkMux
    port map (
            O => \N__50249\,
            I => \N__49819\
        );

    \I__11825\ : ClkMux
    port map (
            O => \N__50248\,
            I => \N__49819\
        );

    \I__11824\ : ClkMux
    port map (
            O => \N__50247\,
            I => \N__49819\
        );

    \I__11823\ : ClkMux
    port map (
            O => \N__50246\,
            I => \N__49819\
        );

    \I__11822\ : ClkMux
    port map (
            O => \N__50245\,
            I => \N__49819\
        );

    \I__11821\ : ClkMux
    port map (
            O => \N__50244\,
            I => \N__49819\
        );

    \I__11820\ : ClkMux
    port map (
            O => \N__50243\,
            I => \N__49819\
        );

    \I__11819\ : ClkMux
    port map (
            O => \N__50242\,
            I => \N__49819\
        );

    \I__11818\ : ClkMux
    port map (
            O => \N__50241\,
            I => \N__49819\
        );

    \I__11817\ : ClkMux
    port map (
            O => \N__50240\,
            I => \N__49819\
        );

    \I__11816\ : ClkMux
    port map (
            O => \N__50239\,
            I => \N__49819\
        );

    \I__11815\ : ClkMux
    port map (
            O => \N__50238\,
            I => \N__49819\
        );

    \I__11814\ : ClkMux
    port map (
            O => \N__50237\,
            I => \N__49819\
        );

    \I__11813\ : ClkMux
    port map (
            O => \N__50236\,
            I => \N__49819\
        );

    \I__11812\ : ClkMux
    port map (
            O => \N__50235\,
            I => \N__49819\
        );

    \I__11811\ : ClkMux
    port map (
            O => \N__50234\,
            I => \N__49819\
        );

    \I__11810\ : ClkMux
    port map (
            O => \N__50233\,
            I => \N__49819\
        );

    \I__11809\ : ClkMux
    port map (
            O => \N__50232\,
            I => \N__49819\
        );

    \I__11808\ : ClkMux
    port map (
            O => \N__50231\,
            I => \N__49819\
        );

    \I__11807\ : ClkMux
    port map (
            O => \N__50230\,
            I => \N__49819\
        );

    \I__11806\ : ClkMux
    port map (
            O => \N__50229\,
            I => \N__49819\
        );

    \I__11805\ : ClkMux
    port map (
            O => \N__50228\,
            I => \N__49819\
        );

    \I__11804\ : ClkMux
    port map (
            O => \N__50227\,
            I => \N__49819\
        );

    \I__11803\ : ClkMux
    port map (
            O => \N__50226\,
            I => \N__49819\
        );

    \I__11802\ : ClkMux
    port map (
            O => \N__50225\,
            I => \N__49819\
        );

    \I__11801\ : ClkMux
    port map (
            O => \N__50224\,
            I => \N__49819\
        );

    \I__11800\ : ClkMux
    port map (
            O => \N__50223\,
            I => \N__49819\
        );

    \I__11799\ : ClkMux
    port map (
            O => \N__50222\,
            I => \N__49819\
        );

    \I__11798\ : ClkMux
    port map (
            O => \N__50221\,
            I => \N__49819\
        );

    \I__11797\ : ClkMux
    port map (
            O => \N__50220\,
            I => \N__49819\
        );

    \I__11796\ : ClkMux
    port map (
            O => \N__50219\,
            I => \N__49819\
        );

    \I__11795\ : ClkMux
    port map (
            O => \N__50218\,
            I => \N__49819\
        );

    \I__11794\ : ClkMux
    port map (
            O => \N__50217\,
            I => \N__49819\
        );

    \I__11793\ : ClkMux
    port map (
            O => \N__50216\,
            I => \N__49819\
        );

    \I__11792\ : ClkMux
    port map (
            O => \N__50215\,
            I => \N__49819\
        );

    \I__11791\ : ClkMux
    port map (
            O => \N__50214\,
            I => \N__49819\
        );

    \I__11790\ : ClkMux
    port map (
            O => \N__50213\,
            I => \N__49819\
        );

    \I__11789\ : ClkMux
    port map (
            O => \N__50212\,
            I => \N__49819\
        );

    \I__11788\ : ClkMux
    port map (
            O => \N__50211\,
            I => \N__49819\
        );

    \I__11787\ : ClkMux
    port map (
            O => \N__50210\,
            I => \N__49819\
        );

    \I__11786\ : ClkMux
    port map (
            O => \N__50209\,
            I => \N__49819\
        );

    \I__11785\ : ClkMux
    port map (
            O => \N__50208\,
            I => \N__49819\
        );

    \I__11784\ : ClkMux
    port map (
            O => \N__50207\,
            I => \N__49819\
        );

    \I__11783\ : ClkMux
    port map (
            O => \N__50206\,
            I => \N__49819\
        );

    \I__11782\ : ClkMux
    port map (
            O => \N__50205\,
            I => \N__49819\
        );

    \I__11781\ : ClkMux
    port map (
            O => \N__50204\,
            I => \N__49819\
        );

    \I__11780\ : ClkMux
    port map (
            O => \N__50203\,
            I => \N__49819\
        );

    \I__11779\ : ClkMux
    port map (
            O => \N__50202\,
            I => \N__49819\
        );

    \I__11778\ : ClkMux
    port map (
            O => \N__50201\,
            I => \N__49819\
        );

    \I__11777\ : ClkMux
    port map (
            O => \N__50200\,
            I => \N__49819\
        );

    \I__11776\ : ClkMux
    port map (
            O => \N__50199\,
            I => \N__49819\
        );

    \I__11775\ : ClkMux
    port map (
            O => \N__50198\,
            I => \N__49819\
        );

    \I__11774\ : ClkMux
    port map (
            O => \N__50197\,
            I => \N__49819\
        );

    \I__11773\ : ClkMux
    port map (
            O => \N__50196\,
            I => \N__49819\
        );

    \I__11772\ : ClkMux
    port map (
            O => \N__50195\,
            I => \N__49819\
        );

    \I__11771\ : ClkMux
    port map (
            O => \N__50194\,
            I => \N__49819\
        );

    \I__11770\ : ClkMux
    port map (
            O => \N__50193\,
            I => \N__49819\
        );

    \I__11769\ : ClkMux
    port map (
            O => \N__50192\,
            I => \N__49819\
        );

    \I__11768\ : ClkMux
    port map (
            O => \N__50191\,
            I => \N__49819\
        );

    \I__11767\ : ClkMux
    port map (
            O => \N__50190\,
            I => \N__49819\
        );

    \I__11766\ : ClkMux
    port map (
            O => \N__50189\,
            I => \N__49819\
        );

    \I__11765\ : ClkMux
    port map (
            O => \N__50188\,
            I => \N__49819\
        );

    \I__11764\ : ClkMux
    port map (
            O => \N__50187\,
            I => \N__49819\
        );

    \I__11763\ : ClkMux
    port map (
            O => \N__50186\,
            I => \N__49819\
        );

    \I__11762\ : ClkMux
    port map (
            O => \N__50185\,
            I => \N__49819\
        );

    \I__11761\ : ClkMux
    port map (
            O => \N__50184\,
            I => \N__49819\
        );

    \I__11760\ : ClkMux
    port map (
            O => \N__50183\,
            I => \N__49819\
        );

    \I__11759\ : ClkMux
    port map (
            O => \N__50182\,
            I => \N__49819\
        );

    \I__11758\ : ClkMux
    port map (
            O => \N__50181\,
            I => \N__49819\
        );

    \I__11757\ : ClkMux
    port map (
            O => \N__50180\,
            I => \N__49819\
        );

    \I__11756\ : ClkMux
    port map (
            O => \N__50179\,
            I => \N__49819\
        );

    \I__11755\ : ClkMux
    port map (
            O => \N__50178\,
            I => \N__49819\
        );

    \I__11754\ : ClkMux
    port map (
            O => \N__50177\,
            I => \N__49819\
        );

    \I__11753\ : ClkMux
    port map (
            O => \N__50176\,
            I => \N__49819\
        );

    \I__11752\ : ClkMux
    port map (
            O => \N__50175\,
            I => \N__49819\
        );

    \I__11751\ : ClkMux
    port map (
            O => \N__50174\,
            I => \N__49819\
        );

    \I__11750\ : ClkMux
    port map (
            O => \N__50173\,
            I => \N__49819\
        );

    \I__11749\ : ClkMux
    port map (
            O => \N__50172\,
            I => \N__49819\
        );

    \I__11748\ : ClkMux
    port map (
            O => \N__50171\,
            I => \N__49819\
        );

    \I__11747\ : ClkMux
    port map (
            O => \N__50170\,
            I => \N__49819\
        );

    \I__11746\ : ClkMux
    port map (
            O => \N__50169\,
            I => \N__49819\
        );

    \I__11745\ : ClkMux
    port map (
            O => \N__50168\,
            I => \N__49819\
        );

    \I__11744\ : ClkMux
    port map (
            O => \N__50167\,
            I => \N__49819\
        );

    \I__11743\ : ClkMux
    port map (
            O => \N__50166\,
            I => \N__49819\
        );

    \I__11742\ : ClkMux
    port map (
            O => \N__50165\,
            I => \N__49819\
        );

    \I__11741\ : ClkMux
    port map (
            O => \N__50164\,
            I => \N__49819\
        );

    \I__11740\ : ClkMux
    port map (
            O => \N__50163\,
            I => \N__49819\
        );

    \I__11739\ : ClkMux
    port map (
            O => \N__50162\,
            I => \N__49819\
        );

    \I__11738\ : ClkMux
    port map (
            O => \N__50161\,
            I => \N__49819\
        );

    \I__11737\ : ClkMux
    port map (
            O => \N__50160\,
            I => \N__49819\
        );

    \I__11736\ : ClkMux
    port map (
            O => \N__50159\,
            I => \N__49819\
        );

    \I__11735\ : ClkMux
    port map (
            O => \N__50158\,
            I => \N__49819\
        );

    \I__11734\ : ClkMux
    port map (
            O => \N__50157\,
            I => \N__49819\
        );

    \I__11733\ : ClkMux
    port map (
            O => \N__50156\,
            I => \N__49819\
        );

    \I__11732\ : ClkMux
    port map (
            O => \N__50155\,
            I => \N__49819\
        );

    \I__11731\ : ClkMux
    port map (
            O => \N__50154\,
            I => \N__49819\
        );

    \I__11730\ : ClkMux
    port map (
            O => \N__50153\,
            I => \N__49819\
        );

    \I__11729\ : ClkMux
    port map (
            O => \N__50152\,
            I => \N__49819\
        );

    \I__11728\ : ClkMux
    port map (
            O => \N__50151\,
            I => \N__49819\
        );

    \I__11727\ : ClkMux
    port map (
            O => \N__50150\,
            I => \N__49819\
        );

    \I__11726\ : ClkMux
    port map (
            O => \N__50149\,
            I => \N__49819\
        );

    \I__11725\ : ClkMux
    port map (
            O => \N__50148\,
            I => \N__49819\
        );

    \I__11724\ : ClkMux
    port map (
            O => \N__50147\,
            I => \N__49819\
        );

    \I__11723\ : ClkMux
    port map (
            O => \N__50146\,
            I => \N__49819\
        );

    \I__11722\ : ClkMux
    port map (
            O => \N__50145\,
            I => \N__49819\
        );

    \I__11721\ : ClkMux
    port map (
            O => \N__50144\,
            I => \N__49819\
        );

    \I__11720\ : ClkMux
    port map (
            O => \N__50143\,
            I => \N__49819\
        );

    \I__11719\ : ClkMux
    port map (
            O => \N__50142\,
            I => \N__49819\
        );

    \I__11718\ : ClkMux
    port map (
            O => \N__50141\,
            I => \N__49819\
        );

    \I__11717\ : ClkMux
    port map (
            O => \N__50140\,
            I => \N__49819\
        );

    \I__11716\ : ClkMux
    port map (
            O => \N__50139\,
            I => \N__49819\
        );

    \I__11715\ : ClkMux
    port map (
            O => \N__50138\,
            I => \N__49819\
        );

    \I__11714\ : ClkMux
    port map (
            O => \N__50137\,
            I => \N__49819\
        );

    \I__11713\ : ClkMux
    port map (
            O => \N__50136\,
            I => \N__49819\
        );

    \I__11712\ : ClkMux
    port map (
            O => \N__50135\,
            I => \N__49819\
        );

    \I__11711\ : ClkMux
    port map (
            O => \N__50134\,
            I => \N__49819\
        );

    \I__11710\ : ClkMux
    port map (
            O => \N__50133\,
            I => \N__49819\
        );

    \I__11709\ : ClkMux
    port map (
            O => \N__50132\,
            I => \N__49819\
        );

    \I__11708\ : ClkMux
    port map (
            O => \N__50131\,
            I => \N__49819\
        );

    \I__11707\ : ClkMux
    port map (
            O => \N__50130\,
            I => \N__49819\
        );

    \I__11706\ : ClkMux
    port map (
            O => \N__50129\,
            I => \N__49819\
        );

    \I__11705\ : ClkMux
    port map (
            O => \N__50128\,
            I => \N__49819\
        );

    \I__11704\ : ClkMux
    port map (
            O => \N__50127\,
            I => \N__49819\
        );

    \I__11703\ : ClkMux
    port map (
            O => \N__50126\,
            I => \N__49819\
        );

    \I__11702\ : GlobalMux
    port map (
            O => \N__49819\,
            I => clk_100mhz_0
        );

    \I__11701\ : CEMux
    port map (
            O => \N__49816\,
            I => \N__49798\
        );

    \I__11700\ : CEMux
    port map (
            O => \N__49815\,
            I => \N__49798\
        );

    \I__11699\ : CEMux
    port map (
            O => \N__49814\,
            I => \N__49798\
        );

    \I__11698\ : CEMux
    port map (
            O => \N__49813\,
            I => \N__49798\
        );

    \I__11697\ : CEMux
    port map (
            O => \N__49812\,
            I => \N__49798\
        );

    \I__11696\ : CEMux
    port map (
            O => \N__49811\,
            I => \N__49798\
        );

    \I__11695\ : GlobalMux
    port map (
            O => \N__49798\,
            I => \N__49795\
        );

    \I__11694\ : gio2CtrlBuf
    port map (
            O => \N__49795\,
            I => \delay_measurement_inst.delay_tr_timer.N_304_i_g\
        );

    \I__11693\ : CascadeMux
    port map (
            O => \N__49792\,
            I => \N__49783\
        );

    \I__11692\ : CascadeMux
    port map (
            O => \N__49791\,
            I => \N__49780\
        );

    \I__11691\ : InMux
    port map (
            O => \N__49790\,
            I => \N__49777\
        );

    \I__11690\ : InMux
    port map (
            O => \N__49789\,
            I => \N__49774\
        );

    \I__11689\ : InMux
    port map (
            O => \N__49788\,
            I => \N__49771\
        );

    \I__11688\ : InMux
    port map (
            O => \N__49787\,
            I => \N__49768\
        );

    \I__11687\ : InMux
    port map (
            O => \N__49786\,
            I => \N__49765\
        );

    \I__11686\ : InMux
    port map (
            O => \N__49783\,
            I => \N__49762\
        );

    \I__11685\ : InMux
    port map (
            O => \N__49780\,
            I => \N__49759\
        );

    \I__11684\ : LocalMux
    port map (
            O => \N__49777\,
            I => \N__49756\
        );

    \I__11683\ : LocalMux
    port map (
            O => \N__49774\,
            I => \N__49753\
        );

    \I__11682\ : LocalMux
    port map (
            O => \N__49771\,
            I => \N__49750\
        );

    \I__11681\ : LocalMux
    port map (
            O => \N__49768\,
            I => \N__49747\
        );

    \I__11680\ : LocalMux
    port map (
            O => \N__49765\,
            I => \N__49657\
        );

    \I__11679\ : LocalMux
    port map (
            O => \N__49762\,
            I => \N__49633\
        );

    \I__11678\ : LocalMux
    port map (
            O => \N__49759\,
            I => \N__49604\
        );

    \I__11677\ : Glb2LocalMux
    port map (
            O => \N__49756\,
            I => \N__49318\
        );

    \I__11676\ : Glb2LocalMux
    port map (
            O => \N__49753\,
            I => \N__49318\
        );

    \I__11675\ : Glb2LocalMux
    port map (
            O => \N__49750\,
            I => \N__49318\
        );

    \I__11674\ : Glb2LocalMux
    port map (
            O => \N__49747\,
            I => \N__49318\
        );

    \I__11673\ : SRMux
    port map (
            O => \N__49746\,
            I => \N__49318\
        );

    \I__11672\ : SRMux
    port map (
            O => \N__49745\,
            I => \N__49318\
        );

    \I__11671\ : SRMux
    port map (
            O => \N__49744\,
            I => \N__49318\
        );

    \I__11670\ : SRMux
    port map (
            O => \N__49743\,
            I => \N__49318\
        );

    \I__11669\ : SRMux
    port map (
            O => \N__49742\,
            I => \N__49318\
        );

    \I__11668\ : SRMux
    port map (
            O => \N__49741\,
            I => \N__49318\
        );

    \I__11667\ : SRMux
    port map (
            O => \N__49740\,
            I => \N__49318\
        );

    \I__11666\ : SRMux
    port map (
            O => \N__49739\,
            I => \N__49318\
        );

    \I__11665\ : SRMux
    port map (
            O => \N__49738\,
            I => \N__49318\
        );

    \I__11664\ : SRMux
    port map (
            O => \N__49737\,
            I => \N__49318\
        );

    \I__11663\ : SRMux
    port map (
            O => \N__49736\,
            I => \N__49318\
        );

    \I__11662\ : SRMux
    port map (
            O => \N__49735\,
            I => \N__49318\
        );

    \I__11661\ : SRMux
    port map (
            O => \N__49734\,
            I => \N__49318\
        );

    \I__11660\ : SRMux
    port map (
            O => \N__49733\,
            I => \N__49318\
        );

    \I__11659\ : SRMux
    port map (
            O => \N__49732\,
            I => \N__49318\
        );

    \I__11658\ : SRMux
    port map (
            O => \N__49731\,
            I => \N__49318\
        );

    \I__11657\ : SRMux
    port map (
            O => \N__49730\,
            I => \N__49318\
        );

    \I__11656\ : SRMux
    port map (
            O => \N__49729\,
            I => \N__49318\
        );

    \I__11655\ : SRMux
    port map (
            O => \N__49728\,
            I => \N__49318\
        );

    \I__11654\ : SRMux
    port map (
            O => \N__49727\,
            I => \N__49318\
        );

    \I__11653\ : SRMux
    port map (
            O => \N__49726\,
            I => \N__49318\
        );

    \I__11652\ : SRMux
    port map (
            O => \N__49725\,
            I => \N__49318\
        );

    \I__11651\ : SRMux
    port map (
            O => \N__49724\,
            I => \N__49318\
        );

    \I__11650\ : SRMux
    port map (
            O => \N__49723\,
            I => \N__49318\
        );

    \I__11649\ : SRMux
    port map (
            O => \N__49722\,
            I => \N__49318\
        );

    \I__11648\ : SRMux
    port map (
            O => \N__49721\,
            I => \N__49318\
        );

    \I__11647\ : SRMux
    port map (
            O => \N__49720\,
            I => \N__49318\
        );

    \I__11646\ : SRMux
    port map (
            O => \N__49719\,
            I => \N__49318\
        );

    \I__11645\ : SRMux
    port map (
            O => \N__49718\,
            I => \N__49318\
        );

    \I__11644\ : SRMux
    port map (
            O => \N__49717\,
            I => \N__49318\
        );

    \I__11643\ : SRMux
    port map (
            O => \N__49716\,
            I => \N__49318\
        );

    \I__11642\ : SRMux
    port map (
            O => \N__49715\,
            I => \N__49318\
        );

    \I__11641\ : SRMux
    port map (
            O => \N__49714\,
            I => \N__49318\
        );

    \I__11640\ : SRMux
    port map (
            O => \N__49713\,
            I => \N__49318\
        );

    \I__11639\ : SRMux
    port map (
            O => \N__49712\,
            I => \N__49318\
        );

    \I__11638\ : SRMux
    port map (
            O => \N__49711\,
            I => \N__49318\
        );

    \I__11637\ : SRMux
    port map (
            O => \N__49710\,
            I => \N__49318\
        );

    \I__11636\ : SRMux
    port map (
            O => \N__49709\,
            I => \N__49318\
        );

    \I__11635\ : SRMux
    port map (
            O => \N__49708\,
            I => \N__49318\
        );

    \I__11634\ : SRMux
    port map (
            O => \N__49707\,
            I => \N__49318\
        );

    \I__11633\ : SRMux
    port map (
            O => \N__49706\,
            I => \N__49318\
        );

    \I__11632\ : SRMux
    port map (
            O => \N__49705\,
            I => \N__49318\
        );

    \I__11631\ : SRMux
    port map (
            O => \N__49704\,
            I => \N__49318\
        );

    \I__11630\ : SRMux
    port map (
            O => \N__49703\,
            I => \N__49318\
        );

    \I__11629\ : SRMux
    port map (
            O => \N__49702\,
            I => \N__49318\
        );

    \I__11628\ : SRMux
    port map (
            O => \N__49701\,
            I => \N__49318\
        );

    \I__11627\ : SRMux
    port map (
            O => \N__49700\,
            I => \N__49318\
        );

    \I__11626\ : SRMux
    port map (
            O => \N__49699\,
            I => \N__49318\
        );

    \I__11625\ : SRMux
    port map (
            O => \N__49698\,
            I => \N__49318\
        );

    \I__11624\ : SRMux
    port map (
            O => \N__49697\,
            I => \N__49318\
        );

    \I__11623\ : SRMux
    port map (
            O => \N__49696\,
            I => \N__49318\
        );

    \I__11622\ : SRMux
    port map (
            O => \N__49695\,
            I => \N__49318\
        );

    \I__11621\ : SRMux
    port map (
            O => \N__49694\,
            I => \N__49318\
        );

    \I__11620\ : SRMux
    port map (
            O => \N__49693\,
            I => \N__49318\
        );

    \I__11619\ : SRMux
    port map (
            O => \N__49692\,
            I => \N__49318\
        );

    \I__11618\ : SRMux
    port map (
            O => \N__49691\,
            I => \N__49318\
        );

    \I__11617\ : SRMux
    port map (
            O => \N__49690\,
            I => \N__49318\
        );

    \I__11616\ : SRMux
    port map (
            O => \N__49689\,
            I => \N__49318\
        );

    \I__11615\ : SRMux
    port map (
            O => \N__49688\,
            I => \N__49318\
        );

    \I__11614\ : SRMux
    port map (
            O => \N__49687\,
            I => \N__49318\
        );

    \I__11613\ : SRMux
    port map (
            O => \N__49686\,
            I => \N__49318\
        );

    \I__11612\ : SRMux
    port map (
            O => \N__49685\,
            I => \N__49318\
        );

    \I__11611\ : SRMux
    port map (
            O => \N__49684\,
            I => \N__49318\
        );

    \I__11610\ : SRMux
    port map (
            O => \N__49683\,
            I => \N__49318\
        );

    \I__11609\ : SRMux
    port map (
            O => \N__49682\,
            I => \N__49318\
        );

    \I__11608\ : SRMux
    port map (
            O => \N__49681\,
            I => \N__49318\
        );

    \I__11607\ : SRMux
    port map (
            O => \N__49680\,
            I => \N__49318\
        );

    \I__11606\ : SRMux
    port map (
            O => \N__49679\,
            I => \N__49318\
        );

    \I__11605\ : SRMux
    port map (
            O => \N__49678\,
            I => \N__49318\
        );

    \I__11604\ : SRMux
    port map (
            O => \N__49677\,
            I => \N__49318\
        );

    \I__11603\ : SRMux
    port map (
            O => \N__49676\,
            I => \N__49318\
        );

    \I__11602\ : SRMux
    port map (
            O => \N__49675\,
            I => \N__49318\
        );

    \I__11601\ : SRMux
    port map (
            O => \N__49674\,
            I => \N__49318\
        );

    \I__11600\ : SRMux
    port map (
            O => \N__49673\,
            I => \N__49318\
        );

    \I__11599\ : SRMux
    port map (
            O => \N__49672\,
            I => \N__49318\
        );

    \I__11598\ : SRMux
    port map (
            O => \N__49671\,
            I => \N__49318\
        );

    \I__11597\ : SRMux
    port map (
            O => \N__49670\,
            I => \N__49318\
        );

    \I__11596\ : SRMux
    port map (
            O => \N__49669\,
            I => \N__49318\
        );

    \I__11595\ : SRMux
    port map (
            O => \N__49668\,
            I => \N__49318\
        );

    \I__11594\ : SRMux
    port map (
            O => \N__49667\,
            I => \N__49318\
        );

    \I__11593\ : SRMux
    port map (
            O => \N__49666\,
            I => \N__49318\
        );

    \I__11592\ : SRMux
    port map (
            O => \N__49665\,
            I => \N__49318\
        );

    \I__11591\ : SRMux
    port map (
            O => \N__49664\,
            I => \N__49318\
        );

    \I__11590\ : SRMux
    port map (
            O => \N__49663\,
            I => \N__49318\
        );

    \I__11589\ : SRMux
    port map (
            O => \N__49662\,
            I => \N__49318\
        );

    \I__11588\ : SRMux
    port map (
            O => \N__49661\,
            I => \N__49318\
        );

    \I__11587\ : SRMux
    port map (
            O => \N__49660\,
            I => \N__49318\
        );

    \I__11586\ : Glb2LocalMux
    port map (
            O => \N__49657\,
            I => \N__49318\
        );

    \I__11585\ : SRMux
    port map (
            O => \N__49656\,
            I => \N__49318\
        );

    \I__11584\ : SRMux
    port map (
            O => \N__49655\,
            I => \N__49318\
        );

    \I__11583\ : SRMux
    port map (
            O => \N__49654\,
            I => \N__49318\
        );

    \I__11582\ : SRMux
    port map (
            O => \N__49653\,
            I => \N__49318\
        );

    \I__11581\ : SRMux
    port map (
            O => \N__49652\,
            I => \N__49318\
        );

    \I__11580\ : SRMux
    port map (
            O => \N__49651\,
            I => \N__49318\
        );

    \I__11579\ : SRMux
    port map (
            O => \N__49650\,
            I => \N__49318\
        );

    \I__11578\ : SRMux
    port map (
            O => \N__49649\,
            I => \N__49318\
        );

    \I__11577\ : SRMux
    port map (
            O => \N__49648\,
            I => \N__49318\
        );

    \I__11576\ : SRMux
    port map (
            O => \N__49647\,
            I => \N__49318\
        );

    \I__11575\ : SRMux
    port map (
            O => \N__49646\,
            I => \N__49318\
        );

    \I__11574\ : SRMux
    port map (
            O => \N__49645\,
            I => \N__49318\
        );

    \I__11573\ : SRMux
    port map (
            O => \N__49644\,
            I => \N__49318\
        );

    \I__11572\ : SRMux
    port map (
            O => \N__49643\,
            I => \N__49318\
        );

    \I__11571\ : SRMux
    port map (
            O => \N__49642\,
            I => \N__49318\
        );

    \I__11570\ : SRMux
    port map (
            O => \N__49641\,
            I => \N__49318\
        );

    \I__11569\ : SRMux
    port map (
            O => \N__49640\,
            I => \N__49318\
        );

    \I__11568\ : SRMux
    port map (
            O => \N__49639\,
            I => \N__49318\
        );

    \I__11567\ : SRMux
    port map (
            O => \N__49638\,
            I => \N__49318\
        );

    \I__11566\ : SRMux
    port map (
            O => \N__49637\,
            I => \N__49318\
        );

    \I__11565\ : SRMux
    port map (
            O => \N__49636\,
            I => \N__49318\
        );

    \I__11564\ : Glb2LocalMux
    port map (
            O => \N__49633\,
            I => \N__49318\
        );

    \I__11563\ : SRMux
    port map (
            O => \N__49632\,
            I => \N__49318\
        );

    \I__11562\ : SRMux
    port map (
            O => \N__49631\,
            I => \N__49318\
        );

    \I__11561\ : SRMux
    port map (
            O => \N__49630\,
            I => \N__49318\
        );

    \I__11560\ : SRMux
    port map (
            O => \N__49629\,
            I => \N__49318\
        );

    \I__11559\ : SRMux
    port map (
            O => \N__49628\,
            I => \N__49318\
        );

    \I__11558\ : SRMux
    port map (
            O => \N__49627\,
            I => \N__49318\
        );

    \I__11557\ : SRMux
    port map (
            O => \N__49626\,
            I => \N__49318\
        );

    \I__11556\ : SRMux
    port map (
            O => \N__49625\,
            I => \N__49318\
        );

    \I__11555\ : SRMux
    port map (
            O => \N__49624\,
            I => \N__49318\
        );

    \I__11554\ : SRMux
    port map (
            O => \N__49623\,
            I => \N__49318\
        );

    \I__11553\ : SRMux
    port map (
            O => \N__49622\,
            I => \N__49318\
        );

    \I__11552\ : SRMux
    port map (
            O => \N__49621\,
            I => \N__49318\
        );

    \I__11551\ : SRMux
    port map (
            O => \N__49620\,
            I => \N__49318\
        );

    \I__11550\ : SRMux
    port map (
            O => \N__49619\,
            I => \N__49318\
        );

    \I__11549\ : SRMux
    port map (
            O => \N__49618\,
            I => \N__49318\
        );

    \I__11548\ : SRMux
    port map (
            O => \N__49617\,
            I => \N__49318\
        );

    \I__11547\ : SRMux
    port map (
            O => \N__49616\,
            I => \N__49318\
        );

    \I__11546\ : SRMux
    port map (
            O => \N__49615\,
            I => \N__49318\
        );

    \I__11545\ : SRMux
    port map (
            O => \N__49614\,
            I => \N__49318\
        );

    \I__11544\ : SRMux
    port map (
            O => \N__49613\,
            I => \N__49318\
        );

    \I__11543\ : SRMux
    port map (
            O => \N__49612\,
            I => \N__49318\
        );

    \I__11542\ : SRMux
    port map (
            O => \N__49611\,
            I => \N__49318\
        );

    \I__11541\ : SRMux
    port map (
            O => \N__49610\,
            I => \N__49318\
        );

    \I__11540\ : SRMux
    port map (
            O => \N__49609\,
            I => \N__49318\
        );

    \I__11539\ : SRMux
    port map (
            O => \N__49608\,
            I => \N__49318\
        );

    \I__11538\ : SRMux
    port map (
            O => \N__49607\,
            I => \N__49318\
        );

    \I__11537\ : Glb2LocalMux
    port map (
            O => \N__49604\,
            I => \N__49318\
        );

    \I__11536\ : SRMux
    port map (
            O => \N__49603\,
            I => \N__49318\
        );

    \I__11535\ : GlobalMux
    port map (
            O => \N__49318\,
            I => \N__49315\
        );

    \I__11534\ : gio2CtrlBuf
    port map (
            O => \N__49315\,
            I => red_c_g
        );

    \I__11533\ : InMux
    port map (
            O => \N__49312\,
            I => \N__49308\
        );

    \I__11532\ : InMux
    port map (
            O => \N__49311\,
            I => \N__49305\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__49308\,
            I => \N__49299\
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__49305\,
            I => \N__49299\
        );

    \I__11529\ : InMux
    port map (
            O => \N__49304\,
            I => \N__49296\
        );

    \I__11528\ : Span4Mux_v
    port map (
            O => \N__49299\,
            I => \N__49293\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__49296\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__11526\ : Odrv4
    port map (
            O => \N__49293\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__11525\ : InMux
    port map (
            O => \N__49288\,
            I => \bfn_18_24_0_\
        );

    \I__11524\ : CascadeMux
    port map (
            O => \N__49285\,
            I => \N__49281\
        );

    \I__11523\ : InMux
    port map (
            O => \N__49284\,
            I => \N__49278\
        );

    \I__11522\ : InMux
    port map (
            O => \N__49281\,
            I => \N__49275\
        );

    \I__11521\ : LocalMux
    port map (
            O => \N__49278\,
            I => \N__49269\
        );

    \I__11520\ : LocalMux
    port map (
            O => \N__49275\,
            I => \N__49269\
        );

    \I__11519\ : InMux
    port map (
            O => \N__49274\,
            I => \N__49266\
        );

    \I__11518\ : Span4Mux_v
    port map (
            O => \N__49269\,
            I => \N__49263\
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__49266\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__11516\ : Odrv4
    port map (
            O => \N__49263\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__11515\ : InMux
    port map (
            O => \N__49258\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__11514\ : CascadeMux
    port map (
            O => \N__49255\,
            I => \N__49251\
        );

    \I__11513\ : CascadeMux
    port map (
            O => \N__49254\,
            I => \N__49248\
        );

    \I__11512\ : InMux
    port map (
            O => \N__49251\,
            I => \N__49243\
        );

    \I__11511\ : InMux
    port map (
            O => \N__49248\,
            I => \N__49243\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__49243\,
            I => \N__49239\
        );

    \I__11509\ : InMux
    port map (
            O => \N__49242\,
            I => \N__49236\
        );

    \I__11508\ : Span4Mux_h
    port map (
            O => \N__49239\,
            I => \N__49233\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__49236\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__11506\ : Odrv4
    port map (
            O => \N__49233\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__11505\ : InMux
    port map (
            O => \N__49228\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__11504\ : CascadeMux
    port map (
            O => \N__49225\,
            I => \N__49221\
        );

    \I__11503\ : CascadeMux
    port map (
            O => \N__49224\,
            I => \N__49218\
        );

    \I__11502\ : InMux
    port map (
            O => \N__49221\,
            I => \N__49213\
        );

    \I__11501\ : InMux
    port map (
            O => \N__49218\,
            I => \N__49213\
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__49213\,
            I => \N__49209\
        );

    \I__11499\ : InMux
    port map (
            O => \N__49212\,
            I => \N__49206\
        );

    \I__11498\ : Span4Mux_h
    port map (
            O => \N__49209\,
            I => \N__49203\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__49206\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__11496\ : Odrv4
    port map (
            O => \N__49203\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__11495\ : InMux
    port map (
            O => \N__49198\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__11494\ : InMux
    port map (
            O => \N__49195\,
            I => \N__49189\
        );

    \I__11493\ : InMux
    port map (
            O => \N__49194\,
            I => \N__49189\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__49189\,
            I => \N__49185\
        );

    \I__11491\ : InMux
    port map (
            O => \N__49188\,
            I => \N__49182\
        );

    \I__11490\ : Span4Mux_h
    port map (
            O => \N__49185\,
            I => \N__49179\
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__49182\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__11488\ : Odrv4
    port map (
            O => \N__49179\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__11487\ : InMux
    port map (
            O => \N__49174\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__11486\ : InMux
    port map (
            O => \N__49171\,
            I => \N__49165\
        );

    \I__11485\ : InMux
    port map (
            O => \N__49170\,
            I => \N__49165\
        );

    \I__11484\ : LocalMux
    port map (
            O => \N__49165\,
            I => \N__49161\
        );

    \I__11483\ : InMux
    port map (
            O => \N__49164\,
            I => \N__49158\
        );

    \I__11482\ : Span4Mux_h
    port map (
            O => \N__49161\,
            I => \N__49155\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__49158\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__11480\ : Odrv4
    port map (
            O => \N__49155\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__11479\ : InMux
    port map (
            O => \N__49150\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__11478\ : CascadeMux
    port map (
            O => \N__49147\,
            I => \N__49143\
        );

    \I__11477\ : CascadeMux
    port map (
            O => \N__49146\,
            I => \N__49140\
        );

    \I__11476\ : InMux
    port map (
            O => \N__49143\,
            I => \N__49134\
        );

    \I__11475\ : InMux
    port map (
            O => \N__49140\,
            I => \N__49134\
        );

    \I__11474\ : InMux
    port map (
            O => \N__49139\,
            I => \N__49131\
        );

    \I__11473\ : LocalMux
    port map (
            O => \N__49134\,
            I => \N__49128\
        );

    \I__11472\ : LocalMux
    port map (
            O => \N__49131\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__11471\ : Odrv12
    port map (
            O => \N__49128\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__11470\ : InMux
    port map (
            O => \N__49123\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__11469\ : CascadeMux
    port map (
            O => \N__49120\,
            I => \N__49116\
        );

    \I__11468\ : CascadeMux
    port map (
            O => \N__49119\,
            I => \N__49113\
        );

    \I__11467\ : InMux
    port map (
            O => \N__49116\,
            I => \N__49107\
        );

    \I__11466\ : InMux
    port map (
            O => \N__49113\,
            I => \N__49107\
        );

    \I__11465\ : InMux
    port map (
            O => \N__49112\,
            I => \N__49104\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__49107\,
            I => \N__49101\
        );

    \I__11463\ : LocalMux
    port map (
            O => \N__49104\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__11462\ : Odrv12
    port map (
            O => \N__49101\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__11461\ : InMux
    port map (
            O => \N__49096\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__11460\ : InMux
    port map (
            O => \N__49093\,
            I => \N__49089\
        );

    \I__11459\ : InMux
    port map (
            O => \N__49092\,
            I => \N__49086\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__49089\,
            I => \N__49080\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__49086\,
            I => \N__49080\
        );

    \I__11456\ : InMux
    port map (
            O => \N__49085\,
            I => \N__49077\
        );

    \I__11455\ : Span4Mux_v
    port map (
            O => \N__49080\,
            I => \N__49074\
        );

    \I__11454\ : LocalMux
    port map (
            O => \N__49077\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__11453\ : Odrv4
    port map (
            O => \N__49074\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__11452\ : InMux
    port map (
            O => \N__49069\,
            I => \bfn_18_25_0_\
        );

    \I__11451\ : CascadeMux
    port map (
            O => \N__49066\,
            I => \N__49062\
        );

    \I__11450\ : InMux
    port map (
            O => \N__49065\,
            I => \N__49058\
        );

    \I__11449\ : InMux
    port map (
            O => \N__49062\,
            I => \N__49055\
        );

    \I__11448\ : InMux
    port map (
            O => \N__49061\,
            I => \N__49052\
        );

    \I__11447\ : LocalMux
    port map (
            O => \N__49058\,
            I => \N__49047\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__49055\,
            I => \N__49047\
        );

    \I__11445\ : LocalMux
    port map (
            O => \N__49052\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__11444\ : Odrv12
    port map (
            O => \N__49047\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__11443\ : InMux
    port map (
            O => \N__49042\,
            I => \bfn_18_23_0_\
        );

    \I__11442\ : InMux
    port map (
            O => \N__49039\,
            I => \N__49034\
        );

    \I__11441\ : InMux
    port map (
            O => \N__49038\,
            I => \N__49031\
        );

    \I__11440\ : InMux
    port map (
            O => \N__49037\,
            I => \N__49028\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__49034\,
            I => \N__49023\
        );

    \I__11438\ : LocalMux
    port map (
            O => \N__49031\,
            I => \N__49023\
        );

    \I__11437\ : LocalMux
    port map (
            O => \N__49028\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__11436\ : Odrv12
    port map (
            O => \N__49023\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__11435\ : InMux
    port map (
            O => \N__49018\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__11434\ : CascadeMux
    port map (
            O => \N__49015\,
            I => \N__49011\
        );

    \I__11433\ : CascadeMux
    port map (
            O => \N__49014\,
            I => \N__49008\
        );

    \I__11432\ : InMux
    port map (
            O => \N__49011\,
            I => \N__49002\
        );

    \I__11431\ : InMux
    port map (
            O => \N__49008\,
            I => \N__49002\
        );

    \I__11430\ : InMux
    port map (
            O => \N__49007\,
            I => \N__48999\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__49002\,
            I => \N__48996\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__48999\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__11427\ : Odrv12
    port map (
            O => \N__48996\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__11426\ : InMux
    port map (
            O => \N__48991\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__11425\ : CascadeMux
    port map (
            O => \N__48988\,
            I => \N__48984\
        );

    \I__11424\ : CascadeMux
    port map (
            O => \N__48987\,
            I => \N__48981\
        );

    \I__11423\ : InMux
    port map (
            O => \N__48984\,
            I => \N__48975\
        );

    \I__11422\ : InMux
    port map (
            O => \N__48981\,
            I => \N__48975\
        );

    \I__11421\ : InMux
    port map (
            O => \N__48980\,
            I => \N__48972\
        );

    \I__11420\ : LocalMux
    port map (
            O => \N__48975\,
            I => \N__48969\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__48972\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__11418\ : Odrv12
    port map (
            O => \N__48969\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__11417\ : InMux
    port map (
            O => \N__48964\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__11416\ : InMux
    port map (
            O => \N__48961\,
            I => \N__48955\
        );

    \I__11415\ : InMux
    port map (
            O => \N__48960\,
            I => \N__48955\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__48955\,
            I => \N__48951\
        );

    \I__11413\ : InMux
    port map (
            O => \N__48954\,
            I => \N__48948\
        );

    \I__11412\ : Span4Mux_h
    port map (
            O => \N__48951\,
            I => \N__48945\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__48948\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__11410\ : Odrv4
    port map (
            O => \N__48945\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__11409\ : InMux
    port map (
            O => \N__48940\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__11408\ : CascadeMux
    port map (
            O => \N__48937\,
            I => \N__48934\
        );

    \I__11407\ : InMux
    port map (
            O => \N__48934\,
            I => \N__48930\
        );

    \I__11406\ : InMux
    port map (
            O => \N__48933\,
            I => \N__48927\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__48930\,
            I => \N__48921\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__48927\,
            I => \N__48921\
        );

    \I__11403\ : InMux
    port map (
            O => \N__48926\,
            I => \N__48918\
        );

    \I__11402\ : Span4Mux_h
    port map (
            O => \N__48921\,
            I => \N__48915\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__48918\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__11400\ : Odrv4
    port map (
            O => \N__48915\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__11399\ : InMux
    port map (
            O => \N__48910\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__11398\ : CascadeMux
    port map (
            O => \N__48907\,
            I => \N__48903\
        );

    \I__11397\ : CascadeMux
    port map (
            O => \N__48906\,
            I => \N__48900\
        );

    \I__11396\ : InMux
    port map (
            O => \N__48903\,
            I => \N__48895\
        );

    \I__11395\ : InMux
    port map (
            O => \N__48900\,
            I => \N__48895\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__48895\,
            I => \N__48891\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48894\,
            I => \N__48888\
        );

    \I__11392\ : Span4Mux_v
    port map (
            O => \N__48891\,
            I => \N__48885\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__48888\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__11390\ : Odrv4
    port map (
            O => \N__48885\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__11389\ : InMux
    port map (
            O => \N__48880\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__11388\ : InMux
    port map (
            O => \N__48877\,
            I => \N__48870\
        );

    \I__11387\ : InMux
    port map (
            O => \N__48876\,
            I => \N__48870\
        );

    \I__11386\ : InMux
    port map (
            O => \N__48875\,
            I => \N__48867\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__48870\,
            I => \N__48864\
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__48867\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__11383\ : Odrv12
    port map (
            O => \N__48864\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__11382\ : InMux
    port map (
            O => \N__48859\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__11381\ : InMux
    port map (
            O => \N__48856\,
            I => \N__48853\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__48853\,
            I => \N__48849\
        );

    \I__11379\ : InMux
    port map (
            O => \N__48852\,
            I => \N__48846\
        );

    \I__11378\ : Span4Mux_h
    port map (
            O => \N__48849\,
            I => \N__48842\
        );

    \I__11377\ : LocalMux
    port map (
            O => \N__48846\,
            I => \N__48839\
        );

    \I__11376\ : InMux
    port map (
            O => \N__48845\,
            I => \N__48836\
        );

    \I__11375\ : Span4Mux_v
    port map (
            O => \N__48842\,
            I => \N__48833\
        );

    \I__11374\ : Span4Mux_h
    port map (
            O => \N__48839\,
            I => \N__48830\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__48836\,
            I => \N__48827\
        );

    \I__11372\ : Span4Mux_h
    port map (
            O => \N__48833\,
            I => \N__48824\
        );

    \I__11371\ : Span4Mux_h
    port map (
            O => \N__48830\,
            I => \N__48819\
        );

    \I__11370\ : Span4Mux_v
    port map (
            O => \N__48827\,
            I => \N__48819\
        );

    \I__11369\ : Odrv4
    port map (
            O => \N__48824\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__11368\ : Odrv4
    port map (
            O => \N__48819\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__11367\ : InMux
    port map (
            O => \N__48814\,
            I => \N__48811\
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__48811\,
            I => \N__48807\
        );

    \I__11365\ : CascadeMux
    port map (
            O => \N__48810\,
            I => \N__48804\
        );

    \I__11364\ : Span4Mux_h
    port map (
            O => \N__48807\,
            I => \N__48801\
        );

    \I__11363\ : InMux
    port map (
            O => \N__48804\,
            I => \N__48798\
        );

    \I__11362\ : Span4Mux_v
    port map (
            O => \N__48801\,
            I => \N__48792\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__48798\,
            I => \N__48792\
        );

    \I__11360\ : InMux
    port map (
            O => \N__48797\,
            I => \N__48789\
        );

    \I__11359\ : Span4Mux_h
    port map (
            O => \N__48792\,
            I => \N__48786\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__48789\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__11357\ : Odrv4
    port map (
            O => \N__48786\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__11356\ : InMux
    port map (
            O => \N__48781\,
            I => \bfn_18_22_0_\
        );

    \I__11355\ : InMux
    port map (
            O => \N__48778\,
            I => \N__48775\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__48775\,
            I => \N__48771\
        );

    \I__11353\ : CascadeMux
    port map (
            O => \N__48774\,
            I => \N__48768\
        );

    \I__11352\ : Span4Mux_h
    port map (
            O => \N__48771\,
            I => \N__48765\
        );

    \I__11351\ : InMux
    port map (
            O => \N__48768\,
            I => \N__48761\
        );

    \I__11350\ : Span4Mux_v
    port map (
            O => \N__48765\,
            I => \N__48758\
        );

    \I__11349\ : InMux
    port map (
            O => \N__48764\,
            I => \N__48755\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__48761\,
            I => \N__48752\
        );

    \I__11347\ : Odrv4
    port map (
            O => \N__48758\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__48755\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__11345\ : Odrv12
    port map (
            O => \N__48752\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__11344\ : InMux
    port map (
            O => \N__48745\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__11343\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48736\
        );

    \I__11342\ : InMux
    port map (
            O => \N__48741\,
            I => \N__48736\
        );

    \I__11341\ : LocalMux
    port map (
            O => \N__48736\,
            I => \N__48732\
        );

    \I__11340\ : InMux
    port map (
            O => \N__48735\,
            I => \N__48729\
        );

    \I__11339\ : Span4Mux_h
    port map (
            O => \N__48732\,
            I => \N__48726\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__48729\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__11337\ : Odrv4
    port map (
            O => \N__48726\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__11336\ : InMux
    port map (
            O => \N__48721\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__11335\ : InMux
    port map (
            O => \N__48718\,
            I => \N__48711\
        );

    \I__11334\ : InMux
    port map (
            O => \N__48717\,
            I => \N__48711\
        );

    \I__11333\ : InMux
    port map (
            O => \N__48716\,
            I => \N__48708\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__48711\,
            I => \N__48705\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__48708\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__11330\ : Odrv12
    port map (
            O => \N__48705\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__11329\ : InMux
    port map (
            O => \N__48700\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__11328\ : CascadeMux
    port map (
            O => \N__48697\,
            I => \N__48693\
        );

    \I__11327\ : CascadeMux
    port map (
            O => \N__48696\,
            I => \N__48690\
        );

    \I__11326\ : InMux
    port map (
            O => \N__48693\,
            I => \N__48684\
        );

    \I__11325\ : InMux
    port map (
            O => \N__48690\,
            I => \N__48684\
        );

    \I__11324\ : InMux
    port map (
            O => \N__48689\,
            I => \N__48681\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__48684\,
            I => \N__48678\
        );

    \I__11322\ : LocalMux
    port map (
            O => \N__48681\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__11321\ : Odrv12
    port map (
            O => \N__48678\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__11320\ : InMux
    port map (
            O => \N__48673\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__11319\ : CascadeMux
    port map (
            O => \N__48670\,
            I => \N__48667\
        );

    \I__11318\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48663\
        );

    \I__11317\ : InMux
    port map (
            O => \N__48666\,
            I => \N__48659\
        );

    \I__11316\ : LocalMux
    port map (
            O => \N__48663\,
            I => \N__48656\
        );

    \I__11315\ : InMux
    port map (
            O => \N__48662\,
            I => \N__48653\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__48659\,
            I => \N__48650\
        );

    \I__11313\ : Span4Mux_h
    port map (
            O => \N__48656\,
            I => \N__48647\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__48653\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__11311\ : Odrv12
    port map (
            O => \N__48650\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__11310\ : Odrv4
    port map (
            O => \N__48647\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__11309\ : InMux
    port map (
            O => \N__48640\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__11308\ : InMux
    port map (
            O => \N__48637\,
            I => \N__48630\
        );

    \I__11307\ : InMux
    port map (
            O => \N__48636\,
            I => \N__48630\
        );

    \I__11306\ : InMux
    port map (
            O => \N__48635\,
            I => \N__48627\
        );

    \I__11305\ : LocalMux
    port map (
            O => \N__48630\,
            I => \N__48624\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__48627\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__11303\ : Odrv12
    port map (
            O => \N__48624\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__11302\ : InMux
    port map (
            O => \N__48619\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__11301\ : CascadeMux
    port map (
            O => \N__48616\,
            I => \N__48612\
        );

    \I__11300\ : CascadeMux
    port map (
            O => \N__48615\,
            I => \N__48609\
        );

    \I__11299\ : InMux
    port map (
            O => \N__48612\,
            I => \N__48604\
        );

    \I__11298\ : InMux
    port map (
            O => \N__48609\,
            I => \N__48604\
        );

    \I__11297\ : LocalMux
    port map (
            O => \N__48604\,
            I => \N__48600\
        );

    \I__11296\ : InMux
    port map (
            O => \N__48603\,
            I => \N__48597\
        );

    \I__11295\ : Span4Mux_v
    port map (
            O => \N__48600\,
            I => \N__48594\
        );

    \I__11294\ : LocalMux
    port map (
            O => \N__48597\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__11293\ : Odrv4
    port map (
            O => \N__48594\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__11292\ : InMux
    port map (
            O => \N__48589\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__11291\ : CascadeMux
    port map (
            O => \N__48586\,
            I => \N__48583\
        );

    \I__11290\ : InMux
    port map (
            O => \N__48583\,
            I => \N__48580\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__48580\,
            I => \N__48575\
        );

    \I__11288\ : InMux
    port map (
            O => \N__48579\,
            I => \N__48572\
        );

    \I__11287\ : InMux
    port map (
            O => \N__48578\,
            I => \N__48569\
        );

    \I__11286\ : Span4Mux_v
    port map (
            O => \N__48575\,
            I => \N__48566\
        );

    \I__11285\ : LocalMux
    port map (
            O => \N__48572\,
            I => \N__48563\
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__48569\,
            I => \N__48560\
        );

    \I__11283\ : Span4Mux_h
    port map (
            O => \N__48566\,
            I => \N__48556\
        );

    \I__11282\ : Span4Mux_v
    port map (
            O => \N__48563\,
            I => \N__48551\
        );

    \I__11281\ : Span4Mux_v
    port map (
            O => \N__48560\,
            I => \N__48551\
        );

    \I__11280\ : InMux
    port map (
            O => \N__48559\,
            I => \N__48548\
        );

    \I__11279\ : Odrv4
    port map (
            O => \N__48556\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__11278\ : Odrv4
    port map (
            O => \N__48551\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__11277\ : LocalMux
    port map (
            O => \N__48548\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__11276\ : InMux
    port map (
            O => \N__48541\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__11275\ : InMux
    port map (
            O => \N__48538\,
            I => \N__48534\
        );

    \I__11274\ : InMux
    port map (
            O => \N__48537\,
            I => \N__48531\
        );

    \I__11273\ : LocalMux
    port map (
            O => \N__48534\,
            I => \N__48524\
        );

    \I__11272\ : LocalMux
    port map (
            O => \N__48531\,
            I => \N__48524\
        );

    \I__11271\ : InMux
    port map (
            O => \N__48530\,
            I => \N__48521\
        );

    \I__11270\ : InMux
    port map (
            O => \N__48529\,
            I => \N__48518\
        );

    \I__11269\ : Span4Mux_v
    port map (
            O => \N__48524\,
            I => \N__48515\
        );

    \I__11268\ : LocalMux
    port map (
            O => \N__48521\,
            I => \N__48512\
        );

    \I__11267\ : LocalMux
    port map (
            O => \N__48518\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__11266\ : Odrv4
    port map (
            O => \N__48515\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__11265\ : Odrv4
    port map (
            O => \N__48512\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__11264\ : InMux
    port map (
            O => \N__48505\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__11263\ : CascadeMux
    port map (
            O => \N__48502\,
            I => \N__48499\
        );

    \I__11262\ : InMux
    port map (
            O => \N__48499\,
            I => \N__48492\
        );

    \I__11261\ : InMux
    port map (
            O => \N__48498\,
            I => \N__48492\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48497\,
            I => \N__48489\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__48492\,
            I => \N__48486\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__48489\,
            I => \N__48482\
        );

    \I__11257\ : Span4Mux_h
    port map (
            O => \N__48486\,
            I => \N__48479\
        );

    \I__11256\ : InMux
    port map (
            O => \N__48485\,
            I => \N__48476\
        );

    \I__11255\ : Odrv12
    port map (
            O => \N__48482\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__11254\ : Odrv4
    port map (
            O => \N__48479\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__11253\ : LocalMux
    port map (
            O => \N__48476\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__11252\ : InMux
    port map (
            O => \N__48469\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__11251\ : InMux
    port map (
            O => \N__48466\,
            I => \N__48462\
        );

    \I__11250\ : InMux
    port map (
            O => \N__48465\,
            I => \N__48459\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__48462\,
            I => \N__48456\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__48459\,
            I => \N__48452\
        );

    \I__11247\ : Span4Mux_h
    port map (
            O => \N__48456\,
            I => \N__48448\
        );

    \I__11246\ : InMux
    port map (
            O => \N__48455\,
            I => \N__48445\
        );

    \I__11245\ : Span4Mux_h
    port map (
            O => \N__48452\,
            I => \N__48442\
        );

    \I__11244\ : InMux
    port map (
            O => \N__48451\,
            I => \N__48439\
        );

    \I__11243\ : Odrv4
    port map (
            O => \N__48448\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__48445\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__11241\ : Odrv4
    port map (
            O => \N__48442\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__11240\ : LocalMux
    port map (
            O => \N__48439\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__11239\ : InMux
    port map (
            O => \N__48430\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__11238\ : InMux
    port map (
            O => \N__48427\,
            I => \N__48423\
        );

    \I__11237\ : InMux
    port map (
            O => \N__48426\,
            I => \N__48420\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__48423\,
            I => \N__48416\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__48420\,
            I => \N__48413\
        );

    \I__11234\ : InMux
    port map (
            O => \N__48419\,
            I => \N__48410\
        );

    \I__11233\ : Span4Mux_v
    port map (
            O => \N__48416\,
            I => \N__48407\
        );

    \I__11232\ : Span4Mux_h
    port map (
            O => \N__48413\,
            I => \N__48404\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__48410\,
            I => \N__48400\
        );

    \I__11230\ : Span4Mux_h
    port map (
            O => \N__48407\,
            I => \N__48395\
        );

    \I__11229\ : Span4Mux_v
    port map (
            O => \N__48404\,
            I => \N__48395\
        );

    \I__11228\ : InMux
    port map (
            O => \N__48403\,
            I => \N__48392\
        );

    \I__11227\ : Odrv4
    port map (
            O => \N__48400\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11226\ : Odrv4
    port map (
            O => \N__48395\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__48392\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11224\ : InMux
    port map (
            O => \N__48385\,
            I => \bfn_18_21_0_\
        );

    \I__11223\ : InMux
    port map (
            O => \N__48382\,
            I => \N__48378\
        );

    \I__11222\ : InMux
    port map (
            O => \N__48381\,
            I => \N__48375\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__48378\,
            I => \N__48370\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__48375\,
            I => \N__48367\
        );

    \I__11219\ : InMux
    port map (
            O => \N__48374\,
            I => \N__48364\
        );

    \I__11218\ : InMux
    port map (
            O => \N__48373\,
            I => \N__48361\
        );

    \I__11217\ : Span4Mux_h
    port map (
            O => \N__48370\,
            I => \N__48356\
        );

    \I__11216\ : Span4Mux_h
    port map (
            O => \N__48367\,
            I => \N__48356\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__48364\,
            I => \N__48353\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__48361\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11213\ : Odrv4
    port map (
            O => \N__48356\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11212\ : Odrv12
    port map (
            O => \N__48353\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11211\ : InMux
    port map (
            O => \N__48346\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__11210\ : InMux
    port map (
            O => \N__48343\,
            I => \N__48338\
        );

    \I__11209\ : InMux
    port map (
            O => \N__48342\,
            I => \N__48333\
        );

    \I__11208\ : InMux
    port map (
            O => \N__48341\,
            I => \N__48333\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__48338\,
            I => \N__48330\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__48333\,
            I => \N__48327\
        );

    \I__11205\ : Span4Mux_h
    port map (
            O => \N__48330\,
            I => \N__48323\
        );

    \I__11204\ : Span4Mux_v
    port map (
            O => \N__48327\,
            I => \N__48320\
        );

    \I__11203\ : InMux
    port map (
            O => \N__48326\,
            I => \N__48317\
        );

    \I__11202\ : Odrv4
    port map (
            O => \N__48323\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__11201\ : Odrv4
    port map (
            O => \N__48320\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__48317\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__11199\ : InMux
    port map (
            O => \N__48310\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__11198\ : InMux
    port map (
            O => \N__48307\,
            I => \N__48304\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__48304\,
            I => \N__48299\
        );

    \I__11196\ : InMux
    port map (
            O => \N__48303\,
            I => \N__48296\
        );

    \I__11195\ : InMux
    port map (
            O => \N__48302\,
            I => \N__48293\
        );

    \I__11194\ : Span4Mux_v
    port map (
            O => \N__48299\,
            I => \N__48288\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__48296\,
            I => \N__48288\
        );

    \I__11192\ : LocalMux
    port map (
            O => \N__48293\,
            I => \N__48285\
        );

    \I__11191\ : Span4Mux_h
    port map (
            O => \N__48288\,
            I => \N__48279\
        );

    \I__11190\ : Span4Mux_v
    port map (
            O => \N__48285\,
            I => \N__48279\
        );

    \I__11189\ : InMux
    port map (
            O => \N__48284\,
            I => \N__48276\
        );

    \I__11188\ : Odrv4
    port map (
            O => \N__48279\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__48276\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__11186\ : InMux
    port map (
            O => \N__48271\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__11185\ : CEMux
    port map (
            O => \N__48268\,
            I => \N__48244\
        );

    \I__11184\ : CEMux
    port map (
            O => \N__48267\,
            I => \N__48244\
        );

    \I__11183\ : CEMux
    port map (
            O => \N__48266\,
            I => \N__48244\
        );

    \I__11182\ : CEMux
    port map (
            O => \N__48265\,
            I => \N__48244\
        );

    \I__11181\ : CEMux
    port map (
            O => \N__48264\,
            I => \N__48244\
        );

    \I__11180\ : CEMux
    port map (
            O => \N__48263\,
            I => \N__48244\
        );

    \I__11179\ : CEMux
    port map (
            O => \N__48262\,
            I => \N__48244\
        );

    \I__11178\ : CEMux
    port map (
            O => \N__48261\,
            I => \N__48244\
        );

    \I__11177\ : GlobalMux
    port map (
            O => \N__48244\,
            I => \N__48241\
        );

    \I__11176\ : gio2CtrlBuf
    port map (
            O => \N__48241\,
            I => \current_shift_inst.timer_s1.N_180_i_g\
        );

    \I__11175\ : InMux
    port map (
            O => \N__48238\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__11174\ : InMux
    port map (
            O => \N__48235\,
            I => \N__48230\
        );

    \I__11173\ : InMux
    port map (
            O => \N__48234\,
            I => \N__48227\
        );

    \I__11172\ : InMux
    port map (
            O => \N__48233\,
            I => \N__48224\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__48230\,
            I => \N__48221\
        );

    \I__11170\ : LocalMux
    port map (
            O => \N__48227\,
            I => \N__48217\
        );

    \I__11169\ : LocalMux
    port map (
            O => \N__48224\,
            I => \N__48214\
        );

    \I__11168\ : Span4Mux_v
    port map (
            O => \N__48221\,
            I => \N__48211\
        );

    \I__11167\ : InMux
    port map (
            O => \N__48220\,
            I => \N__48208\
        );

    \I__11166\ : Span4Mux_v
    port map (
            O => \N__48217\,
            I => \N__48203\
        );

    \I__11165\ : Span4Mux_v
    port map (
            O => \N__48214\,
            I => \N__48203\
        );

    \I__11164\ : Span4Mux_h
    port map (
            O => \N__48211\,
            I => \N__48198\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__48208\,
            I => \N__48198\
        );

    \I__11162\ : Odrv4
    port map (
            O => \N__48203\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__11161\ : Odrv4
    port map (
            O => \N__48198\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__11160\ : InMux
    port map (
            O => \N__48193\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__11159\ : InMux
    port map (
            O => \N__48190\,
            I => \N__48185\
        );

    \I__11158\ : InMux
    port map (
            O => \N__48189\,
            I => \N__48182\
        );

    \I__11157\ : InMux
    port map (
            O => \N__48188\,
            I => \N__48179\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__48185\,
            I => \N__48176\
        );

    \I__11155\ : LocalMux
    port map (
            O => \N__48182\,
            I => \N__48172\
        );

    \I__11154\ : LocalMux
    port map (
            O => \N__48179\,
            I => \N__48169\
        );

    \I__11153\ : Span4Mux_v
    port map (
            O => \N__48176\,
            I => \N__48166\
        );

    \I__11152\ : InMux
    port map (
            O => \N__48175\,
            I => \N__48163\
        );

    \I__11151\ : Span4Mux_v
    port map (
            O => \N__48172\,
            I => \N__48158\
        );

    \I__11150\ : Span4Mux_v
    port map (
            O => \N__48169\,
            I => \N__48158\
        );

    \I__11149\ : Span4Mux_h
    port map (
            O => \N__48166\,
            I => \N__48153\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__48163\,
            I => \N__48153\
        );

    \I__11147\ : Odrv4
    port map (
            O => \N__48158\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__11146\ : Odrv4
    port map (
            O => \N__48153\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__11145\ : InMux
    port map (
            O => \N__48148\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__11144\ : InMux
    port map (
            O => \N__48145\,
            I => \N__48140\
        );

    \I__11143\ : InMux
    port map (
            O => \N__48144\,
            I => \N__48137\
        );

    \I__11142\ : InMux
    port map (
            O => \N__48143\,
            I => \N__48134\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__48140\,
            I => \N__48130\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__48137\,
            I => \N__48127\
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__48134\,
            I => \N__48124\
        );

    \I__11138\ : InMux
    port map (
            O => \N__48133\,
            I => \N__48121\
        );

    \I__11137\ : Span4Mux_h
    port map (
            O => \N__48130\,
            I => \N__48118\
        );

    \I__11136\ : Span4Mux_h
    port map (
            O => \N__48127\,
            I => \N__48115\
        );

    \I__11135\ : Span4Mux_v
    port map (
            O => \N__48124\,
            I => \N__48110\
        );

    \I__11134\ : LocalMux
    port map (
            O => \N__48121\,
            I => \N__48110\
        );

    \I__11133\ : Odrv4
    port map (
            O => \N__48118\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__11132\ : Odrv4
    port map (
            O => \N__48115\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__11131\ : Odrv4
    port map (
            O => \N__48110\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__11130\ : InMux
    port map (
            O => \N__48103\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__11129\ : InMux
    port map (
            O => \N__48100\,
            I => \N__48096\
        );

    \I__11128\ : InMux
    port map (
            O => \N__48099\,
            I => \N__48093\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__48096\,
            I => \N__48090\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__48093\,
            I => \N__48087\
        );

    \I__11125\ : Span4Mux_h
    port map (
            O => \N__48090\,
            I => \N__48082\
        );

    \I__11124\ : Span4Mux_h
    port map (
            O => \N__48087\,
            I => \N__48079\
        );

    \I__11123\ : InMux
    port map (
            O => \N__48086\,
            I => \N__48074\
        );

    \I__11122\ : InMux
    port map (
            O => \N__48085\,
            I => \N__48074\
        );

    \I__11121\ : Odrv4
    port map (
            O => \N__48082\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__11120\ : Odrv4
    port map (
            O => \N__48079\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__11119\ : LocalMux
    port map (
            O => \N__48074\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__11118\ : InMux
    port map (
            O => \N__48067\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__11117\ : CascadeMux
    port map (
            O => \N__48064\,
            I => \N__48061\
        );

    \I__11116\ : InMux
    port map (
            O => \N__48061\,
            I => \N__48058\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__48058\,
            I => \N__48053\
        );

    \I__11114\ : InMux
    port map (
            O => \N__48057\,
            I => \N__48050\
        );

    \I__11113\ : InMux
    port map (
            O => \N__48056\,
            I => \N__48046\
        );

    \I__11112\ : Span4Mux_v
    port map (
            O => \N__48053\,
            I => \N__48043\
        );

    \I__11111\ : LocalMux
    port map (
            O => \N__48050\,
            I => \N__48040\
        );

    \I__11110\ : InMux
    port map (
            O => \N__48049\,
            I => \N__48037\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__48046\,
            I => \N__48034\
        );

    \I__11108\ : Span4Mux_h
    port map (
            O => \N__48043\,
            I => \N__48027\
        );

    \I__11107\ : Span4Mux_v
    port map (
            O => \N__48040\,
            I => \N__48027\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__48037\,
            I => \N__48027\
        );

    \I__11105\ : Odrv4
    port map (
            O => \N__48034\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__11104\ : Odrv4
    port map (
            O => \N__48027\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__11103\ : InMux
    port map (
            O => \N__48022\,
            I => \bfn_18_20_0_\
        );

    \I__11102\ : InMux
    port map (
            O => \N__48019\,
            I => \N__48012\
        );

    \I__11101\ : InMux
    port map (
            O => \N__48018\,
            I => \N__48012\
        );

    \I__11100\ : InMux
    port map (
            O => \N__48017\,
            I => \N__48009\
        );

    \I__11099\ : LocalMux
    port map (
            O => \N__48012\,
            I => \N__48006\
        );

    \I__11098\ : LocalMux
    port map (
            O => \N__48009\,
            I => \N__48002\
        );

    \I__11097\ : Span4Mux_h
    port map (
            O => \N__48006\,
            I => \N__47999\
        );

    \I__11096\ : InMux
    port map (
            O => \N__48005\,
            I => \N__47996\
        );

    \I__11095\ : Odrv4
    port map (
            O => \N__48002\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11094\ : Odrv4
    port map (
            O => \N__47999\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__47996\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11092\ : InMux
    port map (
            O => \N__47989\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__11091\ : CascadeMux
    port map (
            O => \N__47986\,
            I => \N__47982\
        );

    \I__11090\ : InMux
    port map (
            O => \N__47985\,
            I => \N__47978\
        );

    \I__11089\ : InMux
    port map (
            O => \N__47982\,
            I => \N__47973\
        );

    \I__11088\ : InMux
    port map (
            O => \N__47981\,
            I => \N__47973\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__47978\,
            I => \N__47968\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__47973\,
            I => \N__47968\
        );

    \I__11085\ : Span4Mux_v
    port map (
            O => \N__47968\,
            I => \N__47964\
        );

    \I__11084\ : InMux
    port map (
            O => \N__47967\,
            I => \N__47961\
        );

    \I__11083\ : Odrv4
    port map (
            O => \N__47964\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__47961\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__11081\ : InMux
    port map (
            O => \N__47956\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__11080\ : CascadeMux
    port map (
            O => \N__47953\,
            I => \N__47949\
        );

    \I__11079\ : InMux
    port map (
            O => \N__47952\,
            I => \N__47945\
        );

    \I__11078\ : InMux
    port map (
            O => \N__47949\,
            I => \N__47942\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47948\,
            I => \N__47939\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__47945\,
            I => \N__47936\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__47942\,
            I => \N__47933\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__47939\,
            I => \N__47930\
        );

    \I__11073\ : Span4Mux_v
    port map (
            O => \N__47936\,
            I => \N__47927\
        );

    \I__11072\ : Span4Mux_h
    port map (
            O => \N__47933\,
            I => \N__47923\
        );

    \I__11071\ : Span4Mux_v
    port map (
            O => \N__47930\,
            I => \N__47918\
        );

    \I__11070\ : Span4Mux_h
    port map (
            O => \N__47927\,
            I => \N__47918\
        );

    \I__11069\ : InMux
    port map (
            O => \N__47926\,
            I => \N__47915\
        );

    \I__11068\ : Odrv4
    port map (
            O => \N__47923\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__11067\ : Odrv4
    port map (
            O => \N__47918\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__11066\ : LocalMux
    port map (
            O => \N__47915\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__11065\ : InMux
    port map (
            O => \N__47908\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__11064\ : InMux
    port map (
            O => \N__47905\,
            I => \N__47902\
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__47902\,
            I => \N__47897\
        );

    \I__11062\ : InMux
    port map (
            O => \N__47901\,
            I => \N__47894\
        );

    \I__11061\ : InMux
    port map (
            O => \N__47900\,
            I => \N__47890\
        );

    \I__11060\ : Span4Mux_v
    port map (
            O => \N__47897\,
            I => \N__47885\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__47894\,
            I => \N__47885\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47893\,
            I => \N__47882\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__47890\,
            I => \N__47879\
        );

    \I__11056\ : Span4Mux_h
    port map (
            O => \N__47885\,
            I => \N__47876\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__47882\,
            I => \N__47873\
        );

    \I__11054\ : Odrv4
    port map (
            O => \N__47879\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__11053\ : Odrv4
    port map (
            O => \N__47876\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__11052\ : Odrv4
    port map (
            O => \N__47873\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__11051\ : InMux
    port map (
            O => \N__47866\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__11050\ : InMux
    port map (
            O => \N__47863\,
            I => \N__47855\
        );

    \I__11049\ : InMux
    port map (
            O => \N__47862\,
            I => \N__47855\
        );

    \I__11048\ : InMux
    port map (
            O => \N__47861\,
            I => \N__47852\
        );

    \I__11047\ : InMux
    port map (
            O => \N__47860\,
            I => \N__47849\
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__47855\,
            I => \N__47846\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__47852\,
            I => \N__47841\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__47849\,
            I => \N__47841\
        );

    \I__11043\ : Odrv12
    port map (
            O => \N__47846\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__11042\ : Odrv4
    port map (
            O => \N__47841\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__11041\ : InMux
    port map (
            O => \N__47836\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__11040\ : InMux
    port map (
            O => \N__47833\,
            I => \N__47830\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__47830\,
            I => \N__47826\
        );

    \I__11038\ : InMux
    port map (
            O => \N__47829\,
            I => \N__47823\
        );

    \I__11037\ : Span4Mux_v
    port map (
            O => \N__47826\,
            I => \N__47816\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__47823\,
            I => \N__47816\
        );

    \I__11035\ : InMux
    port map (
            O => \N__47822\,
            I => \N__47811\
        );

    \I__11034\ : InMux
    port map (
            O => \N__47821\,
            I => \N__47811\
        );

    \I__11033\ : Span4Mux_h
    port map (
            O => \N__47816\,
            I => \N__47806\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__47811\,
            I => \N__47806\
        );

    \I__11031\ : Odrv4
    port map (
            O => \N__47806\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__11030\ : InMux
    port map (
            O => \N__47803\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__11029\ : InMux
    port map (
            O => \N__47800\,
            I => \N__47797\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__47797\,
            I => \N__47792\
        );

    \I__11027\ : InMux
    port map (
            O => \N__47796\,
            I => \N__47789\
        );

    \I__11026\ : InMux
    port map (
            O => \N__47795\,
            I => \N__47786\
        );

    \I__11025\ : Span4Mux_v
    port map (
            O => \N__47792\,
            I => \N__47780\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__47789\,
            I => \N__47780\
        );

    \I__11023\ : LocalMux
    port map (
            O => \N__47786\,
            I => \N__47777\
        );

    \I__11022\ : InMux
    port map (
            O => \N__47785\,
            I => \N__47774\
        );

    \I__11021\ : Span4Mux_h
    port map (
            O => \N__47780\,
            I => \N__47771\
        );

    \I__11020\ : Span4Mux_h
    port map (
            O => \N__47777\,
            I => \N__47768\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__47774\,
            I => \N__47765\
        );

    \I__11018\ : Odrv4
    port map (
            O => \N__47771\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__11017\ : Odrv4
    port map (
            O => \N__47768\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__11016\ : Odrv12
    port map (
            O => \N__47765\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__11015\ : InMux
    port map (
            O => \N__47758\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__11014\ : InMux
    port map (
            O => \N__47755\,
            I => \N__47752\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__47752\,
            I => \N__47747\
        );

    \I__11012\ : InMux
    port map (
            O => \N__47751\,
            I => \N__47744\
        );

    \I__11011\ : InMux
    port map (
            O => \N__47750\,
            I => \N__47741\
        );

    \I__11010\ : Span4Mux_h
    port map (
            O => \N__47747\,
            I => \N__47736\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__47744\,
            I => \N__47736\
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__47741\,
            I => \N__47733\
        );

    \I__11007\ : Span4Mux_h
    port map (
            O => \N__47736\,
            I => \N__47729\
        );

    \I__11006\ : Span4Mux_h
    port map (
            O => \N__47733\,
            I => \N__47726\
        );

    \I__11005\ : InMux
    port map (
            O => \N__47732\,
            I => \N__47723\
        );

    \I__11004\ : Odrv4
    port map (
            O => \N__47729\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__11003\ : Odrv4
    port map (
            O => \N__47726\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__47723\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__11001\ : InMux
    port map (
            O => \N__47716\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__11000\ : InMux
    port map (
            O => \N__47713\,
            I => \N__47710\
        );

    \I__10999\ : LocalMux
    port map (
            O => \N__47710\,
            I => \N__47705\
        );

    \I__10998\ : InMux
    port map (
            O => \N__47709\,
            I => \N__47702\
        );

    \I__10997\ : InMux
    port map (
            O => \N__47708\,
            I => \N__47698\
        );

    \I__10996\ : Span4Mux_h
    port map (
            O => \N__47705\,
            I => \N__47693\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__47702\,
            I => \N__47693\
        );

    \I__10994\ : InMux
    port map (
            O => \N__47701\,
            I => \N__47690\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__47698\,
            I => \N__47687\
        );

    \I__10992\ : Span4Mux_h
    port map (
            O => \N__47693\,
            I => \N__47682\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__47690\,
            I => \N__47682\
        );

    \I__10990\ : Odrv4
    port map (
            O => \N__47687\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10989\ : Odrv4
    port map (
            O => \N__47682\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10988\ : InMux
    port map (
            O => \N__47677\,
            I => \bfn_18_19_0_\
        );

    \I__10987\ : InMux
    port map (
            O => \N__47674\,
            I => \N__47669\
        );

    \I__10986\ : InMux
    port map (
            O => \N__47673\,
            I => \N__47666\
        );

    \I__10985\ : InMux
    port map (
            O => \N__47672\,
            I => \N__47662\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__47669\,
            I => \N__47659\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__47666\,
            I => \N__47656\
        );

    \I__10982\ : InMux
    port map (
            O => \N__47665\,
            I => \N__47653\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__47662\,
            I => \N__47650\
        );

    \I__10980\ : Span4Mux_v
    port map (
            O => \N__47659\,
            I => \N__47643\
        );

    \I__10979\ : Span4Mux_h
    port map (
            O => \N__47656\,
            I => \N__47643\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__47653\,
            I => \N__47643\
        );

    \I__10977\ : Odrv4
    port map (
            O => \N__47650\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10976\ : Odrv4
    port map (
            O => \N__47643\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10975\ : InMux
    port map (
            O => \N__47638\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__10974\ : CascadeMux
    port map (
            O => \N__47635\,
            I => \N__47632\
        );

    \I__10973\ : InMux
    port map (
            O => \N__47632\,
            I => \N__47627\
        );

    \I__10972\ : InMux
    port map (
            O => \N__47631\,
            I => \N__47624\
        );

    \I__10971\ : InMux
    port map (
            O => \N__47630\,
            I => \N__47621\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__47627\,
            I => \N__47617\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__47624\,
            I => \N__47614\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__47621\,
            I => \N__47611\
        );

    \I__10967\ : InMux
    port map (
            O => \N__47620\,
            I => \N__47608\
        );

    \I__10966\ : Span4Mux_h
    port map (
            O => \N__47617\,
            I => \N__47603\
        );

    \I__10965\ : Span4Mux_v
    port map (
            O => \N__47614\,
            I => \N__47603\
        );

    \I__10964\ : Span4Mux_h
    port map (
            O => \N__47611\,
            I => \N__47598\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__47608\,
            I => \N__47598\
        );

    \I__10962\ : Odrv4
    port map (
            O => \N__47603\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10961\ : Odrv4
    port map (
            O => \N__47598\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10960\ : InMux
    port map (
            O => \N__47593\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__10959\ : InMux
    port map (
            O => \N__47590\,
            I => \N__47587\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__47587\,
            I => \N__47582\
        );

    \I__10957\ : InMux
    port map (
            O => \N__47586\,
            I => \N__47579\
        );

    \I__10956\ : InMux
    port map (
            O => \N__47585\,
            I => \N__47575\
        );

    \I__10955\ : Span4Mux_v
    port map (
            O => \N__47582\,
            I => \N__47570\
        );

    \I__10954\ : LocalMux
    port map (
            O => \N__47579\,
            I => \N__47570\
        );

    \I__10953\ : InMux
    port map (
            O => \N__47578\,
            I => \N__47567\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__47575\,
            I => \N__47564\
        );

    \I__10951\ : Span4Mux_h
    port map (
            O => \N__47570\,
            I => \N__47559\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__47567\,
            I => \N__47559\
        );

    \I__10949\ : Odrv4
    port map (
            O => \N__47564\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10948\ : Odrv4
    port map (
            O => \N__47559\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10947\ : InMux
    port map (
            O => \N__47554\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__10946\ : InMux
    port map (
            O => \N__47551\,
            I => \N__47548\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__47548\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__10944\ : InMux
    port map (
            O => \N__47545\,
            I => \N__47542\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__47542\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__10942\ : InMux
    port map (
            O => \N__47539\,
            I => \N__47536\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__47536\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__10940\ : InMux
    port map (
            O => \N__47533\,
            I => \N__47530\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__47530\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__10938\ : InMux
    port map (
            O => \N__47527\,
            I => \N__47524\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__47524\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__10936\ : CascadeMux
    port map (
            O => \N__47521\,
            I => \N__47518\
        );

    \I__10935\ : InMux
    port map (
            O => \N__47518\,
            I => \N__47512\
        );

    \I__10934\ : InMux
    port map (
            O => \N__47517\,
            I => \N__47512\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__47512\,
            I => \N__47509\
        );

    \I__10932\ : Span4Mux_v
    port map (
            O => \N__47509\,
            I => \N__47504\
        );

    \I__10931\ : InMux
    port map (
            O => \N__47508\,
            I => \N__47501\
        );

    \I__10930\ : InMux
    port map (
            O => \N__47507\,
            I => \N__47498\
        );

    \I__10929\ : Span4Mux_h
    port map (
            O => \N__47504\,
            I => \N__47495\
        );

    \I__10928\ : LocalMux
    port map (
            O => \N__47501\,
            I => \N__47492\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__47498\,
            I => \N__47489\
        );

    \I__10926\ : Odrv4
    port map (
            O => \N__47495\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10925\ : Odrv4
    port map (
            O => \N__47492\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10924\ : Odrv4
    port map (
            O => \N__47489\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10923\ : CascadeMux
    port map (
            O => \N__47482\,
            I => \N__47479\
        );

    \I__10922\ : InMux
    port map (
            O => \N__47479\,
            I => \N__47470\
        );

    \I__10921\ : InMux
    port map (
            O => \N__47478\,
            I => \N__47470\
        );

    \I__10920\ : InMux
    port map (
            O => \N__47477\,
            I => \N__47470\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__47470\,
            I => \N__47466\
        );

    \I__10918\ : InMux
    port map (
            O => \N__47469\,
            I => \N__47463\
        );

    \I__10917\ : Span4Mux_h
    port map (
            O => \N__47466\,
            I => \N__47460\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__47463\,
            I => \N__47457\
        );

    \I__10915\ : Odrv4
    port map (
            O => \N__47460\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__10914\ : Odrv4
    port map (
            O => \N__47457\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__10913\ : InMux
    port map (
            O => \N__47452\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__10912\ : InMux
    port map (
            O => \N__47449\,
            I => \N__47444\
        );

    \I__10911\ : InMux
    port map (
            O => \N__47448\,
            I => \N__47441\
        );

    \I__10910\ : InMux
    port map (
            O => \N__47447\,
            I => \N__47438\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__47444\,
            I => \N__47434\
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__47441\,
            I => \N__47431\
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__47438\,
            I => \N__47428\
        );

    \I__10906\ : InMux
    port map (
            O => \N__47437\,
            I => \N__47425\
        );

    \I__10905\ : Span4Mux_h
    port map (
            O => \N__47434\,
            I => \N__47422\
        );

    \I__10904\ : Span4Mux_v
    port map (
            O => \N__47431\,
            I => \N__47415\
        );

    \I__10903\ : Span4Mux_h
    port map (
            O => \N__47428\,
            I => \N__47415\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__47425\,
            I => \N__47415\
        );

    \I__10901\ : Odrv4
    port map (
            O => \N__47422\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__10900\ : Odrv4
    port map (
            O => \N__47415\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__10899\ : InMux
    port map (
            O => \N__47410\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__10898\ : InMux
    port map (
            O => \N__47407\,
            I => \N__47404\
        );

    \I__10897\ : LocalMux
    port map (
            O => \N__47404\,
            I => \N__47401\
        );

    \I__10896\ : Span4Mux_h
    port map (
            O => \N__47401\,
            I => \N__47396\
        );

    \I__10895\ : InMux
    port map (
            O => \N__47400\,
            I => \N__47393\
        );

    \I__10894\ : InMux
    port map (
            O => \N__47399\,
            I => \N__47390\
        );

    \I__10893\ : Odrv4
    port map (
            O => \N__47396\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__47393\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__47390\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__10890\ : InMux
    port map (
            O => \N__47383\,
            I => \N__47380\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__47380\,
            I => \N__47377\
        );

    \I__10888\ : Span4Mux_v
    port map (
            O => \N__47377\,
            I => \N__47374\
        );

    \I__10887\ : Odrv4
    port map (
            O => \N__47374\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\
        );

    \I__10886\ : CascadeMux
    port map (
            O => \N__47371\,
            I => \N__47368\
        );

    \I__10885\ : InMux
    port map (
            O => \N__47368\,
            I => \N__47365\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__47365\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__10883\ : InMux
    port map (
            O => \N__47362\,
            I => \N__47359\
        );

    \I__10882\ : LocalMux
    port map (
            O => \N__47359\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__10881\ : InMux
    port map (
            O => \N__47356\,
            I => \N__47353\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__47353\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__10879\ : InMux
    port map (
            O => \N__47350\,
            I => \N__47347\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__47347\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__10877\ : InMux
    port map (
            O => \N__47344\,
            I => \N__47341\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__47341\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__10875\ : InMux
    port map (
            O => \N__47338\,
            I => \N__47335\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__47335\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__10873\ : InMux
    port map (
            O => \N__47332\,
            I => \N__47329\
        );

    \I__10872\ : LocalMux
    port map (
            O => \N__47329\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__10871\ : InMux
    port map (
            O => \N__47326\,
            I => \N__47323\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__47323\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__10869\ : InMux
    port map (
            O => \N__47320\,
            I => \N__47317\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__47317\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__10867\ : InMux
    port map (
            O => \N__47314\,
            I => \N__47308\
        );

    \I__10866\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47308\
        );

    \I__10865\ : LocalMux
    port map (
            O => \N__47308\,
            I => \N__47305\
        );

    \I__10864\ : Span4Mux_h
    port map (
            O => \N__47305\,
            I => \N__47302\
        );

    \I__10863\ : Span4Mux_h
    port map (
            O => \N__47302\,
            I => \N__47297\
        );

    \I__10862\ : InMux
    port map (
            O => \N__47301\,
            I => \N__47292\
        );

    \I__10861\ : InMux
    port map (
            O => \N__47300\,
            I => \N__47292\
        );

    \I__10860\ : Odrv4
    port map (
            O => \N__47297\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__47292\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10858\ : InMux
    port map (
            O => \N__47287\,
            I => \N__47284\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__47284\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__10856\ : InMux
    port map (
            O => \N__47281\,
            I => \N__47254\
        );

    \I__10855\ : InMux
    port map (
            O => \N__47280\,
            I => \N__47254\
        );

    \I__10854\ : InMux
    port map (
            O => \N__47279\,
            I => \N__47254\
        );

    \I__10853\ : InMux
    port map (
            O => \N__47278\,
            I => \N__47254\
        );

    \I__10852\ : InMux
    port map (
            O => \N__47277\,
            I => \N__47254\
        );

    \I__10851\ : InMux
    port map (
            O => \N__47276\,
            I => \N__47251\
        );

    \I__10850\ : InMux
    port map (
            O => \N__47275\,
            I => \N__47246\
        );

    \I__10849\ : InMux
    port map (
            O => \N__47274\,
            I => \N__47246\
        );

    \I__10848\ : InMux
    port map (
            O => \N__47273\,
            I => \N__47241\
        );

    \I__10847\ : InMux
    port map (
            O => \N__47272\,
            I => \N__47241\
        );

    \I__10846\ : InMux
    port map (
            O => \N__47271\,
            I => \N__47234\
        );

    \I__10845\ : InMux
    port map (
            O => \N__47270\,
            I => \N__47234\
        );

    \I__10844\ : InMux
    port map (
            O => \N__47269\,
            I => \N__47234\
        );

    \I__10843\ : InMux
    port map (
            O => \N__47268\,
            I => \N__47227\
        );

    \I__10842\ : InMux
    port map (
            O => \N__47267\,
            I => \N__47227\
        );

    \I__10841\ : InMux
    port map (
            O => \N__47266\,
            I => \N__47227\
        );

    \I__10840\ : InMux
    port map (
            O => \N__47265\,
            I => \N__47220\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__47254\,
            I => \N__47216\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__47251\,
            I => \N__47212\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__47246\,
            I => \N__47203\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__47241\,
            I => \N__47203\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__47234\,
            I => \N__47203\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__47227\,
            I => \N__47203\
        );

    \I__10833\ : InMux
    port map (
            O => \N__47226\,
            I => \N__47198\
        );

    \I__10832\ : InMux
    port map (
            O => \N__47225\,
            I => \N__47198\
        );

    \I__10831\ : InMux
    port map (
            O => \N__47224\,
            I => \N__47193\
        );

    \I__10830\ : InMux
    port map (
            O => \N__47223\,
            I => \N__47193\
        );

    \I__10829\ : LocalMux
    port map (
            O => \N__47220\,
            I => \N__47189\
        );

    \I__10828\ : InMux
    port map (
            O => \N__47219\,
            I => \N__47185\
        );

    \I__10827\ : Span4Mux_h
    port map (
            O => \N__47216\,
            I => \N__47182\
        );

    \I__10826\ : InMux
    port map (
            O => \N__47215\,
            I => \N__47179\
        );

    \I__10825\ : Span4Mux_v
    port map (
            O => \N__47212\,
            I => \N__47170\
        );

    \I__10824\ : Span4Mux_v
    port map (
            O => \N__47203\,
            I => \N__47170\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__47198\,
            I => \N__47170\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__47193\,
            I => \N__47170\
        );

    \I__10821\ : InMux
    port map (
            O => \N__47192\,
            I => \N__47167\
        );

    \I__10820\ : Span4Mux_h
    port map (
            O => \N__47189\,
            I => \N__47164\
        );

    \I__10819\ : InMux
    port map (
            O => \N__47188\,
            I => \N__47161\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__47185\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10817\ : Odrv4
    port map (
            O => \N__47182\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__47179\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10815\ : Odrv4
    port map (
            O => \N__47170\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__47167\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10813\ : Odrv4
    port map (
            O => \N__47164\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__47161\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10811\ : InMux
    port map (
            O => \N__47146\,
            I => \N__47140\
        );

    \I__10810\ : InMux
    port map (
            O => \N__47145\,
            I => \N__47140\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__47140\,
            I => \N__47137\
        );

    \I__10808\ : Span12Mux_v
    port map (
            O => \N__47137\,
            I => \N__47133\
        );

    \I__10807\ : InMux
    port map (
            O => \N__47136\,
            I => \N__47130\
        );

    \I__10806\ : Odrv12
    port map (
            O => \N__47133\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__47130\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__10804\ : InMux
    port map (
            O => \N__47125\,
            I => \N__47122\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__47122\,
            I => \N__47119\
        );

    \I__10802\ : Odrv4
    port map (
            O => \N__47119\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__10801\ : InMux
    port map (
            O => \N__47116\,
            I => \N__47113\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__47113\,
            I => \N__47108\
        );

    \I__10799\ : InMux
    port map (
            O => \N__47112\,
            I => \N__47105\
        );

    \I__10798\ : InMux
    port map (
            O => \N__47111\,
            I => \N__47102\
        );

    \I__10797\ : Odrv4
    port map (
            O => \N__47108\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__47105\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__47102\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10794\ : InMux
    port map (
            O => \N__47095\,
            I => \N__47092\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__47092\,
            I => \N__47089\
        );

    \I__10792\ : Span4Mux_h
    port map (
            O => \N__47089\,
            I => \N__47086\
        );

    \I__10791\ : Span4Mux_h
    port map (
            O => \N__47086\,
            I => \N__47083\
        );

    \I__10790\ : Odrv4
    port map (
            O => \N__47083\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\
        );

    \I__10789\ : InMux
    port map (
            O => \N__47080\,
            I => \N__47073\
        );

    \I__10788\ : InMux
    port map (
            O => \N__47079\,
            I => \N__47073\
        );

    \I__10787\ : InMux
    port map (
            O => \N__47078\,
            I => \N__47070\
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__47073\,
            I => \N__47067\
        );

    \I__10785\ : LocalMux
    port map (
            O => \N__47070\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__10784\ : Odrv4
    port map (
            O => \N__47067\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__10783\ : InMux
    port map (
            O => \N__47062\,
            I => \N__47059\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__47059\,
            I => \N__47056\
        );

    \I__10781\ : Span4Mux_v
    port map (
            O => \N__47056\,
            I => \N__47053\
        );

    \I__10780\ : Odrv4
    port map (
            O => \N__47053\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\
        );

    \I__10779\ : InMux
    port map (
            O => \N__47050\,
            I => \N__47047\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__47047\,
            I => \N__47044\
        );

    \I__10777\ : Span4Mux_h
    port map (
            O => \N__47044\,
            I => \N__47041\
        );

    \I__10776\ : Span4Mux_h
    port map (
            O => \N__47041\,
            I => \N__47038\
        );

    \I__10775\ : Odrv4
    port map (
            O => \N__47038\,
            I => \current_shift_inst.un38_control_input_0_s0_11\
        );

    \I__10774\ : InMux
    port map (
            O => \N__47035\,
            I => \N__47032\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__47032\,
            I => \N__47029\
        );

    \I__10772\ : Span4Mux_h
    port map (
            O => \N__47029\,
            I => \N__47026\
        );

    \I__10771\ : Span4Mux_v
    port map (
            O => \N__47026\,
            I => \N__47023\
        );

    \I__10770\ : Odrv4
    port map (
            O => \N__47023\,
            I => \current_shift_inst.un38_control_input_0_s1_11\
        );

    \I__10769\ : InMux
    port map (
            O => \N__47020\,
            I => \N__47017\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__47017\,
            I => \N__47014\
        );

    \I__10767\ : Odrv12
    port map (
            O => \N__47014\,
            I => \current_shift_inst.control_input_1_axb_5\
        );

    \I__10766\ : InMux
    port map (
            O => \N__47011\,
            I => \N__47008\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__47008\,
            I => \N__47005\
        );

    \I__10764\ : Span4Mux_v
    port map (
            O => \N__47005\,
            I => \N__47002\
        );

    \I__10763\ : Span4Mux_h
    port map (
            O => \N__47002\,
            I => \N__46999\
        );

    \I__10762\ : Odrv4
    port map (
            O => \N__46999\,
            I => \current_shift_inst.un38_control_input_0_s0_13\
        );

    \I__10761\ : CascadeMux
    port map (
            O => \N__46996\,
            I => \N__46988\
        );

    \I__10760\ : InMux
    port map (
            O => \N__46995\,
            I => \N__46981\
        );

    \I__10759\ : InMux
    port map (
            O => \N__46994\,
            I => \N__46981\
        );

    \I__10758\ : InMux
    port map (
            O => \N__46993\,
            I => \N__46981\
        );

    \I__10757\ : CascadeMux
    port map (
            O => \N__46992\,
            I => \N__46976\
        );

    \I__10756\ : CascadeMux
    port map (
            O => \N__46991\,
            I => \N__46966\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46988\,
            I => \N__46962\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__46981\,
            I => \N__46959\
        );

    \I__10753\ : InMux
    port map (
            O => \N__46980\,
            I => \N__46950\
        );

    \I__10752\ : InMux
    port map (
            O => \N__46979\,
            I => \N__46950\
        );

    \I__10751\ : InMux
    port map (
            O => \N__46976\,
            I => \N__46950\
        );

    \I__10750\ : InMux
    port map (
            O => \N__46975\,
            I => \N__46950\
        );

    \I__10749\ : InMux
    port map (
            O => \N__46974\,
            I => \N__46937\
        );

    \I__10748\ : InMux
    port map (
            O => \N__46973\,
            I => \N__46937\
        );

    \I__10747\ : InMux
    port map (
            O => \N__46972\,
            I => \N__46937\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46971\,
            I => \N__46937\
        );

    \I__10745\ : InMux
    port map (
            O => \N__46970\,
            I => \N__46937\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46969\,
            I => \N__46937\
        );

    \I__10743\ : InMux
    port map (
            O => \N__46966\,
            I => \N__46932\
        );

    \I__10742\ : InMux
    port map (
            O => \N__46965\,
            I => \N__46932\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__46962\,
            I => \N__46921\
        );

    \I__10740\ : Span4Mux_h
    port map (
            O => \N__46959\,
            I => \N__46918\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__46950\,
            I => \N__46915\
        );

    \I__10738\ : LocalMux
    port map (
            O => \N__46937\,
            I => \N__46912\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__46932\,
            I => \N__46909\
        );

    \I__10736\ : CascadeMux
    port map (
            O => \N__46931\,
            I => \N__46906\
        );

    \I__10735\ : CascadeMux
    port map (
            O => \N__46930\,
            I => \N__46903\
        );

    \I__10734\ : CascadeMux
    port map (
            O => \N__46929\,
            I => \N__46898\
        );

    \I__10733\ : InMux
    port map (
            O => \N__46928\,
            I => \N__46886\
        );

    \I__10732\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46886\
        );

    \I__10731\ : InMux
    port map (
            O => \N__46926\,
            I => \N__46886\
        );

    \I__10730\ : InMux
    port map (
            O => \N__46925\,
            I => \N__46886\
        );

    \I__10729\ : InMux
    port map (
            O => \N__46924\,
            I => \N__46886\
        );

    \I__10728\ : Span4Mux_v
    port map (
            O => \N__46921\,
            I => \N__46881\
        );

    \I__10727\ : Span4Mux_v
    port map (
            O => \N__46918\,
            I => \N__46881\
        );

    \I__10726\ : Span4Mux_h
    port map (
            O => \N__46915\,
            I => \N__46878\
        );

    \I__10725\ : Span4Mux_h
    port map (
            O => \N__46912\,
            I => \N__46873\
        );

    \I__10724\ : Span4Mux_h
    port map (
            O => \N__46909\,
            I => \N__46873\
        );

    \I__10723\ : InMux
    port map (
            O => \N__46906\,
            I => \N__46860\
        );

    \I__10722\ : InMux
    port map (
            O => \N__46903\,
            I => \N__46860\
        );

    \I__10721\ : InMux
    port map (
            O => \N__46902\,
            I => \N__46860\
        );

    \I__10720\ : InMux
    port map (
            O => \N__46901\,
            I => \N__46860\
        );

    \I__10719\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46860\
        );

    \I__10718\ : InMux
    port map (
            O => \N__46897\,
            I => \N__46860\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__46886\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10716\ : Odrv4
    port map (
            O => \N__46881\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10715\ : Odrv4
    port map (
            O => \N__46878\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10714\ : Odrv4
    port map (
            O => \N__46873\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10713\ : LocalMux
    port map (
            O => \N__46860\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10712\ : InMux
    port map (
            O => \N__46849\,
            I => \N__46846\
        );

    \I__10711\ : LocalMux
    port map (
            O => \N__46846\,
            I => \N__46843\
        );

    \I__10710\ : Span4Mux_h
    port map (
            O => \N__46843\,
            I => \N__46840\
        );

    \I__10709\ : Span4Mux_v
    port map (
            O => \N__46840\,
            I => \N__46837\
        );

    \I__10708\ : Odrv4
    port map (
            O => \N__46837\,
            I => \current_shift_inst.un38_control_input_0_s1_13\
        );

    \I__10707\ : InMux
    port map (
            O => \N__46834\,
            I => \N__46831\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__46831\,
            I => \N__46828\
        );

    \I__10705\ : Odrv12
    port map (
            O => \N__46828\,
            I => \current_shift_inst.control_input_1_axb_7\
        );

    \I__10704\ : InMux
    port map (
            O => \N__46825\,
            I => \N__46822\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__46822\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__10702\ : InMux
    port map (
            O => \N__46819\,
            I => \N__46804\
        );

    \I__10701\ : InMux
    port map (
            O => \N__46818\,
            I => \N__46804\
        );

    \I__10700\ : InMux
    port map (
            O => \N__46817\,
            I => \N__46791\
        );

    \I__10699\ : InMux
    port map (
            O => \N__46816\,
            I => \N__46791\
        );

    \I__10698\ : InMux
    port map (
            O => \N__46815\,
            I => \N__46788\
        );

    \I__10697\ : InMux
    port map (
            O => \N__46814\,
            I => \N__46785\
        );

    \I__10696\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46774\
        );

    \I__10695\ : InMux
    port map (
            O => \N__46812\,
            I => \N__46774\
        );

    \I__10694\ : InMux
    port map (
            O => \N__46811\,
            I => \N__46774\
        );

    \I__10693\ : InMux
    port map (
            O => \N__46810\,
            I => \N__46774\
        );

    \I__10692\ : InMux
    port map (
            O => \N__46809\,
            I => \N__46774\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__46804\,
            I => \N__46768\
        );

    \I__10690\ : InMux
    port map (
            O => \N__46803\,
            I => \N__46765\
        );

    \I__10689\ : InMux
    port map (
            O => \N__46802\,
            I => \N__46762\
        );

    \I__10688\ : InMux
    port map (
            O => \N__46801\,
            I => \N__46759\
        );

    \I__10687\ : InMux
    port map (
            O => \N__46800\,
            I => \N__46753\
        );

    \I__10686\ : InMux
    port map (
            O => \N__46799\,
            I => \N__46750\
        );

    \I__10685\ : InMux
    port map (
            O => \N__46798\,
            I => \N__46746\
        );

    \I__10684\ : CascadeMux
    port map (
            O => \N__46797\,
            I => \N__46736\
        );

    \I__10683\ : InMux
    port map (
            O => \N__46796\,
            I => \N__46733\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__46791\,
            I => \N__46724\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__46788\,
            I => \N__46724\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__46785\,
            I => \N__46724\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__46774\,
            I => \N__46724\
        );

    \I__10678\ : InMux
    port map (
            O => \N__46773\,
            I => \N__46717\
        );

    \I__10677\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46717\
        );

    \I__10676\ : InMux
    port map (
            O => \N__46771\,
            I => \N__46717\
        );

    \I__10675\ : Span4Mux_v
    port map (
            O => \N__46768\,
            I => \N__46708\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__46765\,
            I => \N__46708\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__46762\,
            I => \N__46708\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__46759\,
            I => \N__46708\
        );

    \I__10671\ : InMux
    port map (
            O => \N__46758\,
            I => \N__46671\
        );

    \I__10670\ : InMux
    port map (
            O => \N__46757\,
            I => \N__46671\
        );

    \I__10669\ : InMux
    port map (
            O => \N__46756\,
            I => \N__46671\
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__46753\,
            I => \N__46668\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__46750\,
            I => \N__46665\
        );

    \I__10666\ : InMux
    port map (
            O => \N__46749\,
            I => \N__46662\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__46746\,
            I => \N__46659\
        );

    \I__10664\ : InMux
    port map (
            O => \N__46745\,
            I => \N__46652\
        );

    \I__10663\ : InMux
    port map (
            O => \N__46744\,
            I => \N__46652\
        );

    \I__10662\ : InMux
    port map (
            O => \N__46743\,
            I => \N__46652\
        );

    \I__10661\ : CascadeMux
    port map (
            O => \N__46742\,
            I => \N__46648\
        );

    \I__10660\ : InMux
    port map (
            O => \N__46741\,
            I => \N__46644\
        );

    \I__10659\ : InMux
    port map (
            O => \N__46740\,
            I => \N__46639\
        );

    \I__10658\ : InMux
    port map (
            O => \N__46739\,
            I => \N__46639\
        );

    \I__10657\ : InMux
    port map (
            O => \N__46736\,
            I => \N__46636\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__46733\,
            I => \N__46633\
        );

    \I__10655\ : Span4Mux_v
    port map (
            O => \N__46724\,
            I => \N__46628\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__46717\,
            I => \N__46628\
        );

    \I__10653\ : Span4Mux_v
    port map (
            O => \N__46708\,
            I => \N__46625\
        );

    \I__10652\ : InMux
    port map (
            O => \N__46707\,
            I => \N__46622\
        );

    \I__10651\ : InMux
    port map (
            O => \N__46706\,
            I => \N__46617\
        );

    \I__10650\ : InMux
    port map (
            O => \N__46705\,
            I => \N__46617\
        );

    \I__10649\ : InMux
    port map (
            O => \N__46704\,
            I => \N__46614\
        );

    \I__10648\ : InMux
    port map (
            O => \N__46703\,
            I => \N__46609\
        );

    \I__10647\ : InMux
    port map (
            O => \N__46702\,
            I => \N__46609\
        );

    \I__10646\ : InMux
    port map (
            O => \N__46701\,
            I => \N__46604\
        );

    \I__10645\ : InMux
    port map (
            O => \N__46700\,
            I => \N__46604\
        );

    \I__10644\ : InMux
    port map (
            O => \N__46699\,
            I => \N__46593\
        );

    \I__10643\ : InMux
    port map (
            O => \N__46698\,
            I => \N__46593\
        );

    \I__10642\ : InMux
    port map (
            O => \N__46697\,
            I => \N__46593\
        );

    \I__10641\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46593\
        );

    \I__10640\ : InMux
    port map (
            O => \N__46695\,
            I => \N__46593\
        );

    \I__10639\ : InMux
    port map (
            O => \N__46694\,
            I => \N__46586\
        );

    \I__10638\ : InMux
    port map (
            O => \N__46693\,
            I => \N__46586\
        );

    \I__10637\ : InMux
    port map (
            O => \N__46692\,
            I => \N__46586\
        );

    \I__10636\ : InMux
    port map (
            O => \N__46691\,
            I => \N__46577\
        );

    \I__10635\ : InMux
    port map (
            O => \N__46690\,
            I => \N__46577\
        );

    \I__10634\ : InMux
    port map (
            O => \N__46689\,
            I => \N__46577\
        );

    \I__10633\ : InMux
    port map (
            O => \N__46688\,
            I => \N__46577\
        );

    \I__10632\ : InMux
    port map (
            O => \N__46687\,
            I => \N__46566\
        );

    \I__10631\ : InMux
    port map (
            O => \N__46686\,
            I => \N__46566\
        );

    \I__10630\ : InMux
    port map (
            O => \N__46685\,
            I => \N__46566\
        );

    \I__10629\ : InMux
    port map (
            O => \N__46684\,
            I => \N__46566\
        );

    \I__10628\ : InMux
    port map (
            O => \N__46683\,
            I => \N__46566\
        );

    \I__10627\ : InMux
    port map (
            O => \N__46682\,
            I => \N__46561\
        );

    \I__10626\ : InMux
    port map (
            O => \N__46681\,
            I => \N__46561\
        );

    \I__10625\ : InMux
    port map (
            O => \N__46680\,
            I => \N__46554\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46679\,
            I => \N__46554\
        );

    \I__10623\ : InMux
    port map (
            O => \N__46678\,
            I => \N__46554\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__46671\,
            I => \N__46551\
        );

    \I__10621\ : Span4Mux_v
    port map (
            O => \N__46668\,
            I => \N__46544\
        );

    \I__10620\ : Span4Mux_h
    port map (
            O => \N__46665\,
            I => \N__46544\
        );

    \I__10619\ : LocalMux
    port map (
            O => \N__46662\,
            I => \N__46544\
        );

    \I__10618\ : Span4Mux_h
    port map (
            O => \N__46659\,
            I => \N__46539\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__46652\,
            I => \N__46539\
        );

    \I__10616\ : InMux
    port map (
            O => \N__46651\,
            I => \N__46532\
        );

    \I__10615\ : InMux
    port map (
            O => \N__46648\,
            I => \N__46532\
        );

    \I__10614\ : InMux
    port map (
            O => \N__46647\,
            I => \N__46532\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__46644\,
            I => \N__46522\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__46639\,
            I => \N__46522\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__46636\,
            I => \N__46517\
        );

    \I__10610\ : Span4Mux_h
    port map (
            O => \N__46633\,
            I => \N__46517\
        );

    \I__10609\ : Span4Mux_h
    port map (
            O => \N__46628\,
            I => \N__46514\
        );

    \I__10608\ : Sp12to4
    port map (
            O => \N__46625\,
            I => \N__46507\
        );

    \I__10607\ : LocalMux
    port map (
            O => \N__46622\,
            I => \N__46507\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__46617\,
            I => \N__46507\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__46614\,
            I => \N__46504\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__46609\,
            I => \N__46501\
        );

    \I__10603\ : LocalMux
    port map (
            O => \N__46604\,
            I => \N__46490\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__46593\,
            I => \N__46490\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__46586\,
            I => \N__46490\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__46577\,
            I => \N__46490\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__46566\,
            I => \N__46490\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__46561\,
            I => \N__46485\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__46554\,
            I => \N__46485\
        );

    \I__10596\ : Span4Mux_h
    port map (
            O => \N__46551\,
            I => \N__46482\
        );

    \I__10595\ : Span4Mux_h
    port map (
            O => \N__46544\,
            I => \N__46477\
        );

    \I__10594\ : Span4Mux_h
    port map (
            O => \N__46539\,
            I => \N__46477\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__46532\,
            I => \N__46474\
        );

    \I__10592\ : InMux
    port map (
            O => \N__46531\,
            I => \N__46467\
        );

    \I__10591\ : InMux
    port map (
            O => \N__46530\,
            I => \N__46467\
        );

    \I__10590\ : InMux
    port map (
            O => \N__46529\,
            I => \N__46467\
        );

    \I__10589\ : InMux
    port map (
            O => \N__46528\,
            I => \N__46462\
        );

    \I__10588\ : InMux
    port map (
            O => \N__46527\,
            I => \N__46462\
        );

    \I__10587\ : Span4Mux_h
    port map (
            O => \N__46522\,
            I => \N__46457\
        );

    \I__10586\ : Span4Mux_h
    port map (
            O => \N__46517\,
            I => \N__46457\
        );

    \I__10585\ : Sp12to4
    port map (
            O => \N__46514\,
            I => \N__46452\
        );

    \I__10584\ : Span12Mux_h
    port map (
            O => \N__46507\,
            I => \N__46452\
        );

    \I__10583\ : Span4Mux_h
    port map (
            O => \N__46504\,
            I => \N__46443\
        );

    \I__10582\ : Span4Mux_h
    port map (
            O => \N__46501\,
            I => \N__46443\
        );

    \I__10581\ : Span4Mux_v
    port map (
            O => \N__46490\,
            I => \N__46443\
        );

    \I__10580\ : Span4Mux_v
    port map (
            O => \N__46485\,
            I => \N__46443\
        );

    \I__10579\ : Span4Mux_h
    port map (
            O => \N__46482\,
            I => \N__46440\
        );

    \I__10578\ : Odrv4
    port map (
            O => \N__46477\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10577\ : Odrv4
    port map (
            O => \N__46474\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__46467\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__46462\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10574\ : Odrv4
    port map (
            O => \N__46457\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10573\ : Odrv12
    port map (
            O => \N__46452\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10572\ : Odrv4
    port map (
            O => \N__46443\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10571\ : Odrv4
    port map (
            O => \N__46440\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10570\ : CascadeMux
    port map (
            O => \N__46423\,
            I => \N__46415\
        );

    \I__10569\ : CascadeMux
    port map (
            O => \N__46422\,
            I => \N__46412\
        );

    \I__10568\ : CascadeMux
    port map (
            O => \N__46421\,
            I => \N__46409\
        );

    \I__10567\ : CascadeMux
    port map (
            O => \N__46420\,
            I => \N__46403\
        );

    \I__10566\ : CascadeMux
    port map (
            O => \N__46419\,
            I => \N__46400\
        );

    \I__10565\ : CascadeMux
    port map (
            O => \N__46418\,
            I => \N__46397\
        );

    \I__10564\ : InMux
    port map (
            O => \N__46415\,
            I => \N__46392\
        );

    \I__10563\ : InMux
    port map (
            O => \N__46412\,
            I => \N__46392\
        );

    \I__10562\ : InMux
    port map (
            O => \N__46409\,
            I => \N__46389\
        );

    \I__10561\ : CascadeMux
    port map (
            O => \N__46408\,
            I => \N__46386\
        );

    \I__10560\ : CascadeMux
    port map (
            O => \N__46407\,
            I => \N__46383\
        );

    \I__10559\ : CascadeMux
    port map (
            O => \N__46406\,
            I => \N__46380\
        );

    \I__10558\ : InMux
    port map (
            O => \N__46403\,
            I => \N__46363\
        );

    \I__10557\ : InMux
    port map (
            O => \N__46400\,
            I => \N__46358\
        );

    \I__10556\ : InMux
    port map (
            O => \N__46397\,
            I => \N__46358\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__46392\,
            I => \N__46353\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__46389\,
            I => \N__46353\
        );

    \I__10553\ : InMux
    port map (
            O => \N__46386\,
            I => \N__46348\
        );

    \I__10552\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46348\
        );

    \I__10551\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46345\
        );

    \I__10550\ : CascadeMux
    port map (
            O => \N__46379\,
            I => \N__46336\
        );

    \I__10549\ : CascadeMux
    port map (
            O => \N__46378\,
            I => \N__46316\
        );

    \I__10548\ : CascadeMux
    port map (
            O => \N__46377\,
            I => \N__46312\
        );

    \I__10547\ : CascadeMux
    port map (
            O => \N__46376\,
            I => \N__46309\
        );

    \I__10546\ : CascadeMux
    port map (
            O => \N__46375\,
            I => \N__46306\
        );

    \I__10545\ : CascadeMux
    port map (
            O => \N__46374\,
            I => \N__46298\
        );

    \I__10544\ : CascadeMux
    port map (
            O => \N__46373\,
            I => \N__46287\
        );

    \I__10543\ : CascadeMux
    port map (
            O => \N__46372\,
            I => \N__46284\
        );

    \I__10542\ : CascadeMux
    port map (
            O => \N__46371\,
            I => \N__46280\
        );

    \I__10541\ : CascadeMux
    port map (
            O => \N__46370\,
            I => \N__46277\
        );

    \I__10540\ : CascadeMux
    port map (
            O => \N__46369\,
            I => \N__46270\
        );

    \I__10539\ : CascadeMux
    port map (
            O => \N__46368\,
            I => \N__46267\
        );

    \I__10538\ : CascadeMux
    port map (
            O => \N__46367\,
            I => \N__46264\
        );

    \I__10537\ : CascadeMux
    port map (
            O => \N__46366\,
            I => \N__46261\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__46363\,
            I => \N__46250\
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__46358\,
            I => \N__46250\
        );

    \I__10534\ : Span4Mux_h
    port map (
            O => \N__46353\,
            I => \N__46243\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__46348\,
            I => \N__46243\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__46345\,
            I => \N__46243\
        );

    \I__10531\ : CascadeMux
    port map (
            O => \N__46344\,
            I => \N__46240\
        );

    \I__10530\ : CascadeMux
    port map (
            O => \N__46343\,
            I => \N__46237\
        );

    \I__10529\ : CascadeMux
    port map (
            O => \N__46342\,
            I => \N__46234\
        );

    \I__10528\ : CascadeMux
    port map (
            O => \N__46341\,
            I => \N__46225\
        );

    \I__10527\ : CascadeMux
    port map (
            O => \N__46340\,
            I => \N__46222\
        );

    \I__10526\ : InMux
    port map (
            O => \N__46339\,
            I => \N__46219\
        );

    \I__10525\ : InMux
    port map (
            O => \N__46336\,
            I => \N__46205\
        );

    \I__10524\ : CascadeMux
    port map (
            O => \N__46335\,
            I => \N__46202\
        );

    \I__10523\ : CascadeMux
    port map (
            O => \N__46334\,
            I => \N__46199\
        );

    \I__10522\ : CascadeMux
    port map (
            O => \N__46333\,
            I => \N__46196\
        );

    \I__10521\ : CascadeMux
    port map (
            O => \N__46332\,
            I => \N__46193\
        );

    \I__10520\ : CascadeMux
    port map (
            O => \N__46331\,
            I => \N__46190\
        );

    \I__10519\ : CascadeMux
    port map (
            O => \N__46330\,
            I => \N__46187\
        );

    \I__10518\ : CascadeMux
    port map (
            O => \N__46329\,
            I => \N__46184\
        );

    \I__10517\ : CascadeMux
    port map (
            O => \N__46328\,
            I => \N__46181\
        );

    \I__10516\ : CascadeMux
    port map (
            O => \N__46327\,
            I => \N__46178\
        );

    \I__10515\ : CascadeMux
    port map (
            O => \N__46326\,
            I => \N__46175\
        );

    \I__10514\ : CascadeMux
    port map (
            O => \N__46325\,
            I => \N__46172\
        );

    \I__10513\ : CascadeMux
    port map (
            O => \N__46324\,
            I => \N__46169\
        );

    \I__10512\ : CascadeMux
    port map (
            O => \N__46323\,
            I => \N__46165\
        );

    \I__10511\ : CascadeMux
    port map (
            O => \N__46322\,
            I => \N__46162\
        );

    \I__10510\ : CascadeMux
    port map (
            O => \N__46321\,
            I => \N__46159\
        );

    \I__10509\ : CascadeMux
    port map (
            O => \N__46320\,
            I => \N__46156\
        );

    \I__10508\ : CascadeMux
    port map (
            O => \N__46319\,
            I => \N__46153\
        );

    \I__10507\ : InMux
    port map (
            O => \N__46316\,
            I => \N__46149\
        );

    \I__10506\ : InMux
    port map (
            O => \N__46315\,
            I => \N__46140\
        );

    \I__10505\ : InMux
    port map (
            O => \N__46312\,
            I => \N__46140\
        );

    \I__10504\ : InMux
    port map (
            O => \N__46309\,
            I => \N__46140\
        );

    \I__10503\ : InMux
    port map (
            O => \N__46306\,
            I => \N__46140\
        );

    \I__10502\ : CascadeMux
    port map (
            O => \N__46305\,
            I => \N__46137\
        );

    \I__10501\ : CascadeMux
    port map (
            O => \N__46304\,
            I => \N__46134\
        );

    \I__10500\ : CascadeMux
    port map (
            O => \N__46303\,
            I => \N__46131\
        );

    \I__10499\ : CascadeMux
    port map (
            O => \N__46302\,
            I => \N__46128\
        );

    \I__10498\ : InMux
    port map (
            O => \N__46301\,
            I => \N__46123\
        );

    \I__10497\ : InMux
    port map (
            O => \N__46298\,
            I => \N__46123\
        );

    \I__10496\ : CascadeMux
    port map (
            O => \N__46297\,
            I => \N__46120\
        );

    \I__10495\ : CascadeMux
    port map (
            O => \N__46296\,
            I => \N__46117\
        );

    \I__10494\ : CascadeMux
    port map (
            O => \N__46295\,
            I => \N__46114\
        );

    \I__10493\ : CascadeMux
    port map (
            O => \N__46294\,
            I => \N__46111\
        );

    \I__10492\ : CascadeMux
    port map (
            O => \N__46293\,
            I => \N__46108\
        );

    \I__10491\ : CascadeMux
    port map (
            O => \N__46292\,
            I => \N__46105\
        );

    \I__10490\ : CascadeMux
    port map (
            O => \N__46291\,
            I => \N__46102\
        );

    \I__10489\ : CascadeMux
    port map (
            O => \N__46290\,
            I => \N__46099\
        );

    \I__10488\ : InMux
    port map (
            O => \N__46287\,
            I => \N__46095\
        );

    \I__10487\ : InMux
    port map (
            O => \N__46284\,
            I => \N__46086\
        );

    \I__10486\ : InMux
    port map (
            O => \N__46283\,
            I => \N__46086\
        );

    \I__10485\ : InMux
    port map (
            O => \N__46280\,
            I => \N__46086\
        );

    \I__10484\ : InMux
    port map (
            O => \N__46277\,
            I => \N__46086\
        );

    \I__10483\ : CascadeMux
    port map (
            O => \N__46276\,
            I => \N__46083\
        );

    \I__10482\ : CascadeMux
    port map (
            O => \N__46275\,
            I => \N__46080\
        );

    \I__10481\ : CascadeMux
    port map (
            O => \N__46274\,
            I => \N__46077\
        );

    \I__10480\ : CascadeMux
    port map (
            O => \N__46273\,
            I => \N__46074\
        );

    \I__10479\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46065\
        );

    \I__10478\ : InMux
    port map (
            O => \N__46267\,
            I => \N__46065\
        );

    \I__10477\ : InMux
    port map (
            O => \N__46264\,
            I => \N__46065\
        );

    \I__10476\ : InMux
    port map (
            O => \N__46261\,
            I => \N__46065\
        );

    \I__10475\ : CascadeMux
    port map (
            O => \N__46260\,
            I => \N__46062\
        );

    \I__10474\ : CascadeMux
    port map (
            O => \N__46259\,
            I => \N__46059\
        );

    \I__10473\ : CascadeMux
    port map (
            O => \N__46258\,
            I => \N__46056\
        );

    \I__10472\ : CascadeMux
    port map (
            O => \N__46257\,
            I => \N__46053\
        );

    \I__10471\ : CascadeMux
    port map (
            O => \N__46256\,
            I => \N__46050\
        );

    \I__10470\ : CascadeMux
    port map (
            O => \N__46255\,
            I => \N__46047\
        );

    \I__10469\ : Span4Mux_v
    port map (
            O => \N__46250\,
            I => \N__46042\
        );

    \I__10468\ : Span4Mux_v
    port map (
            O => \N__46243\,
            I => \N__46042\
        );

    \I__10467\ : InMux
    port map (
            O => \N__46240\,
            I => \N__46039\
        );

    \I__10466\ : InMux
    port map (
            O => \N__46237\,
            I => \N__46034\
        );

    \I__10465\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46034\
        );

    \I__10464\ : InMux
    port map (
            O => \N__46233\,
            I => \N__46027\
        );

    \I__10463\ : InMux
    port map (
            O => \N__46232\,
            I => \N__46027\
        );

    \I__10462\ : InMux
    port map (
            O => \N__46231\,
            I => \N__46027\
        );

    \I__10461\ : CascadeMux
    port map (
            O => \N__46230\,
            I => \N__46023\
        );

    \I__10460\ : CascadeMux
    port map (
            O => \N__46229\,
            I => \N__46020\
        );

    \I__10459\ : CascadeMux
    port map (
            O => \N__46228\,
            I => \N__46016\
        );

    \I__10458\ : InMux
    port map (
            O => \N__46225\,
            I => \N__46011\
        );

    \I__10457\ : InMux
    port map (
            O => \N__46222\,
            I => \N__46011\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__46219\,
            I => \N__46008\
        );

    \I__10455\ : CascadeMux
    port map (
            O => \N__46218\,
            I => \N__46003\
        );

    \I__10454\ : CascadeMux
    port map (
            O => \N__46217\,
            I => \N__46000\
        );

    \I__10453\ : CascadeMux
    port map (
            O => \N__46216\,
            I => \N__45988\
        );

    \I__10452\ : CascadeMux
    port map (
            O => \N__46215\,
            I => \N__45985\
        );

    \I__10451\ : CascadeMux
    port map (
            O => \N__46214\,
            I => \N__45982\
        );

    \I__10450\ : CascadeMux
    port map (
            O => \N__46213\,
            I => \N__45978\
        );

    \I__10449\ : CascadeMux
    port map (
            O => \N__46212\,
            I => \N__45975\
        );

    \I__10448\ : CascadeMux
    port map (
            O => \N__46211\,
            I => \N__45972\
        );

    \I__10447\ : CascadeMux
    port map (
            O => \N__46210\,
            I => \N__45968\
        );

    \I__10446\ : CascadeMux
    port map (
            O => \N__46209\,
            I => \N__45964\
        );

    \I__10445\ : CascadeMux
    port map (
            O => \N__46208\,
            I => \N__45960\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__46205\,
            I => \N__45956\
        );

    \I__10443\ : InMux
    port map (
            O => \N__46202\,
            I => \N__45949\
        );

    \I__10442\ : InMux
    port map (
            O => \N__46199\,
            I => \N__45949\
        );

    \I__10441\ : InMux
    port map (
            O => \N__46196\,
            I => \N__45949\
        );

    \I__10440\ : InMux
    port map (
            O => \N__46193\,
            I => \N__45940\
        );

    \I__10439\ : InMux
    port map (
            O => \N__46190\,
            I => \N__45940\
        );

    \I__10438\ : InMux
    port map (
            O => \N__46187\,
            I => \N__45940\
        );

    \I__10437\ : InMux
    port map (
            O => \N__46184\,
            I => \N__45940\
        );

    \I__10436\ : InMux
    port map (
            O => \N__46181\,
            I => \N__45931\
        );

    \I__10435\ : InMux
    port map (
            O => \N__46178\,
            I => \N__45931\
        );

    \I__10434\ : InMux
    port map (
            O => \N__46175\,
            I => \N__45931\
        );

    \I__10433\ : InMux
    port map (
            O => \N__46172\,
            I => \N__45931\
        );

    \I__10432\ : InMux
    port map (
            O => \N__46169\,
            I => \N__45922\
        );

    \I__10431\ : CascadeMux
    port map (
            O => \N__46168\,
            I => \N__45918\
        );

    \I__10430\ : InMux
    port map (
            O => \N__46165\,
            I => \N__45913\
        );

    \I__10429\ : InMux
    port map (
            O => \N__46162\,
            I => \N__45913\
        );

    \I__10428\ : InMux
    port map (
            O => \N__46159\,
            I => \N__45906\
        );

    \I__10427\ : InMux
    port map (
            O => \N__46156\,
            I => \N__45906\
        );

    \I__10426\ : InMux
    port map (
            O => \N__46153\,
            I => \N__45906\
        );

    \I__10425\ : InMux
    port map (
            O => \N__46152\,
            I => \N__45903\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__46149\,
            I => \N__45898\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__46140\,
            I => \N__45898\
        );

    \I__10422\ : InMux
    port map (
            O => \N__46137\,
            I => \N__45889\
        );

    \I__10421\ : InMux
    port map (
            O => \N__46134\,
            I => \N__45889\
        );

    \I__10420\ : InMux
    port map (
            O => \N__46131\,
            I => \N__45889\
        );

    \I__10419\ : InMux
    port map (
            O => \N__46128\,
            I => \N__45889\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__46123\,
            I => \N__45886\
        );

    \I__10417\ : InMux
    port map (
            O => \N__46120\,
            I => \N__45877\
        );

    \I__10416\ : InMux
    port map (
            O => \N__46117\,
            I => \N__45877\
        );

    \I__10415\ : InMux
    port map (
            O => \N__46114\,
            I => \N__45877\
        );

    \I__10414\ : InMux
    port map (
            O => \N__46111\,
            I => \N__45877\
        );

    \I__10413\ : InMux
    port map (
            O => \N__46108\,
            I => \N__45870\
        );

    \I__10412\ : InMux
    port map (
            O => \N__46105\,
            I => \N__45870\
        );

    \I__10411\ : InMux
    port map (
            O => \N__46102\,
            I => \N__45870\
        );

    \I__10410\ : InMux
    port map (
            O => \N__46099\,
            I => \N__45865\
        );

    \I__10409\ : InMux
    port map (
            O => \N__46098\,
            I => \N__45865\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__46095\,
            I => \N__45860\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__46086\,
            I => \N__45860\
        );

    \I__10406\ : InMux
    port map (
            O => \N__46083\,
            I => \N__45851\
        );

    \I__10405\ : InMux
    port map (
            O => \N__46080\,
            I => \N__45851\
        );

    \I__10404\ : InMux
    port map (
            O => \N__46077\,
            I => \N__45851\
        );

    \I__10403\ : InMux
    port map (
            O => \N__46074\,
            I => \N__45851\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__46065\,
            I => \N__45848\
        );

    \I__10401\ : InMux
    port map (
            O => \N__46062\,
            I => \N__45841\
        );

    \I__10400\ : InMux
    port map (
            O => \N__46059\,
            I => \N__45841\
        );

    \I__10399\ : InMux
    port map (
            O => \N__46056\,
            I => \N__45841\
        );

    \I__10398\ : InMux
    port map (
            O => \N__46053\,
            I => \N__45834\
        );

    \I__10397\ : InMux
    port map (
            O => \N__46050\,
            I => \N__45834\
        );

    \I__10396\ : InMux
    port map (
            O => \N__46047\,
            I => \N__45834\
        );

    \I__10395\ : Span4Mux_h
    port map (
            O => \N__46042\,
            I => \N__45825\
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__46039\,
            I => \N__45825\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__46034\,
            I => \N__45825\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__46027\,
            I => \N__45825\
        );

    \I__10391\ : InMux
    port map (
            O => \N__46026\,
            I => \N__45822\
        );

    \I__10390\ : InMux
    port map (
            O => \N__46023\,
            I => \N__45817\
        );

    \I__10389\ : InMux
    port map (
            O => \N__46020\,
            I => \N__45817\
        );

    \I__10388\ : CascadeMux
    port map (
            O => \N__46019\,
            I => \N__45814\
        );

    \I__10387\ : InMux
    port map (
            O => \N__46016\,
            I => \N__45811\
        );

    \I__10386\ : LocalMux
    port map (
            O => \N__46011\,
            I => \N__45806\
        );

    \I__10385\ : Span4Mux_h
    port map (
            O => \N__46008\,
            I => \N__45806\
        );

    \I__10384\ : InMux
    port map (
            O => \N__46007\,
            I => \N__45801\
        );

    \I__10383\ : InMux
    port map (
            O => \N__46006\,
            I => \N__45801\
        );

    \I__10382\ : InMux
    port map (
            O => \N__46003\,
            I => \N__45796\
        );

    \I__10381\ : InMux
    port map (
            O => \N__46000\,
            I => \N__45796\
        );

    \I__10380\ : InMux
    port map (
            O => \N__45999\,
            I => \N__45793\
        );

    \I__10379\ : CascadeMux
    port map (
            O => \N__45998\,
            I => \N__45790\
        );

    \I__10378\ : CascadeMux
    port map (
            O => \N__45997\,
            I => \N__45787\
        );

    \I__10377\ : CascadeMux
    port map (
            O => \N__45996\,
            I => \N__45784\
        );

    \I__10376\ : CascadeMux
    port map (
            O => \N__45995\,
            I => \N__45781\
        );

    \I__10375\ : CascadeMux
    port map (
            O => \N__45994\,
            I => \N__45778\
        );

    \I__10374\ : CascadeMux
    port map (
            O => \N__45993\,
            I => \N__45775\
        );

    \I__10373\ : CascadeMux
    port map (
            O => \N__45992\,
            I => \N__45772\
        );

    \I__10372\ : CascadeMux
    port map (
            O => \N__45991\,
            I => \N__45769\
        );

    \I__10371\ : InMux
    port map (
            O => \N__45988\,
            I => \N__45764\
        );

    \I__10370\ : InMux
    port map (
            O => \N__45985\,
            I => \N__45764\
        );

    \I__10369\ : InMux
    port map (
            O => \N__45982\,
            I => \N__45753\
        );

    \I__10368\ : InMux
    port map (
            O => \N__45981\,
            I => \N__45753\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45978\,
            I => \N__45753\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45975\,
            I => \N__45753\
        );

    \I__10365\ : InMux
    port map (
            O => \N__45972\,
            I => \N__45753\
        );

    \I__10364\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45738\
        );

    \I__10363\ : InMux
    port map (
            O => \N__45968\,
            I => \N__45738\
        );

    \I__10362\ : InMux
    port map (
            O => \N__45967\,
            I => \N__45738\
        );

    \I__10361\ : InMux
    port map (
            O => \N__45964\,
            I => \N__45738\
        );

    \I__10360\ : InMux
    port map (
            O => \N__45963\,
            I => \N__45738\
        );

    \I__10359\ : InMux
    port map (
            O => \N__45960\,
            I => \N__45738\
        );

    \I__10358\ : InMux
    port map (
            O => \N__45959\,
            I => \N__45738\
        );

    \I__10357\ : Span4Mux_h
    port map (
            O => \N__45956\,
            I => \N__45729\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__45949\,
            I => \N__45729\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__45940\,
            I => \N__45729\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__45931\,
            I => \N__45729\
        );

    \I__10353\ : CascadeMux
    port map (
            O => \N__45930\,
            I => \N__45726\
        );

    \I__10352\ : CascadeMux
    port map (
            O => \N__45929\,
            I => \N__45723\
        );

    \I__10351\ : CascadeMux
    port map (
            O => \N__45928\,
            I => \N__45720\
        );

    \I__10350\ : CascadeMux
    port map (
            O => \N__45927\,
            I => \N__45717\
        );

    \I__10349\ : CascadeMux
    port map (
            O => \N__45926\,
            I => \N__45714\
        );

    \I__10348\ : CascadeMux
    port map (
            O => \N__45925\,
            I => \N__45711\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__45922\,
            I => \N__45708\
        );

    \I__10346\ : InMux
    port map (
            O => \N__45921\,
            I => \N__45703\
        );

    \I__10345\ : InMux
    port map (
            O => \N__45918\,
            I => \N__45703\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__45913\,
            I => \N__45694\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__45906\,
            I => \N__45694\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__45903\,
            I => \N__45694\
        );

    \I__10341\ : Span4Mux_v
    port map (
            O => \N__45898\,
            I => \N__45694\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__45889\,
            I => \N__45673\
        );

    \I__10339\ : Span4Mux_v
    port map (
            O => \N__45886\,
            I => \N__45673\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__45877\,
            I => \N__45673\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__45870\,
            I => \N__45673\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__45865\,
            I => \N__45673\
        );

    \I__10335\ : Span4Mux_v
    port map (
            O => \N__45860\,
            I => \N__45673\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__45851\,
            I => \N__45673\
        );

    \I__10333\ : Span4Mux_h
    port map (
            O => \N__45848\,
            I => \N__45673\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__45841\,
            I => \N__45673\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__45834\,
            I => \N__45673\
        );

    \I__10330\ : Span4Mux_v
    port map (
            O => \N__45825\,
            I => \N__45670\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__45822\,
            I => \N__45667\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__45817\,
            I => \N__45664\
        );

    \I__10327\ : InMux
    port map (
            O => \N__45814\,
            I => \N__45661\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__45811\,
            I => \N__45656\
        );

    \I__10325\ : Span4Mux_h
    port map (
            O => \N__45806\,
            I => \N__45656\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__45801\,
            I => \N__45649\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__45796\,
            I => \N__45649\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__45793\,
            I => \N__45649\
        );

    \I__10321\ : InMux
    port map (
            O => \N__45790\,
            I => \N__45640\
        );

    \I__10320\ : InMux
    port map (
            O => \N__45787\,
            I => \N__45640\
        );

    \I__10319\ : InMux
    port map (
            O => \N__45784\,
            I => \N__45640\
        );

    \I__10318\ : InMux
    port map (
            O => \N__45781\,
            I => \N__45640\
        );

    \I__10317\ : InMux
    port map (
            O => \N__45778\,
            I => \N__45631\
        );

    \I__10316\ : InMux
    port map (
            O => \N__45775\,
            I => \N__45631\
        );

    \I__10315\ : InMux
    port map (
            O => \N__45772\,
            I => \N__45631\
        );

    \I__10314\ : InMux
    port map (
            O => \N__45769\,
            I => \N__45631\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__45764\,
            I => \N__45622\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__45753\,
            I => \N__45622\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__45738\,
            I => \N__45622\
        );

    \I__10310\ : Span4Mux_h
    port map (
            O => \N__45729\,
            I => \N__45622\
        );

    \I__10309\ : InMux
    port map (
            O => \N__45726\,
            I => \N__45615\
        );

    \I__10308\ : InMux
    port map (
            O => \N__45723\,
            I => \N__45615\
        );

    \I__10307\ : InMux
    port map (
            O => \N__45720\,
            I => \N__45615\
        );

    \I__10306\ : InMux
    port map (
            O => \N__45717\,
            I => \N__45608\
        );

    \I__10305\ : InMux
    port map (
            O => \N__45714\,
            I => \N__45608\
        );

    \I__10304\ : InMux
    port map (
            O => \N__45711\,
            I => \N__45608\
        );

    \I__10303\ : Span4Mux_h
    port map (
            O => \N__45708\,
            I => \N__45599\
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__45703\,
            I => \N__45599\
        );

    \I__10301\ : Span4Mux_v
    port map (
            O => \N__45694\,
            I => \N__45599\
        );

    \I__10300\ : Span4Mux_v
    port map (
            O => \N__45673\,
            I => \N__45599\
        );

    \I__10299\ : Odrv4
    port map (
            O => \N__45670\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10298\ : Odrv12
    port map (
            O => \N__45667\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10297\ : Odrv12
    port map (
            O => \N__45664\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__45661\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10295\ : Odrv4
    port map (
            O => \N__45656\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10294\ : Odrv12
    port map (
            O => \N__45649\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__45640\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__45631\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10291\ : Odrv4
    port map (
            O => \N__45622\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__45615\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__45608\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__45599\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10287\ : InMux
    port map (
            O => \N__45574\,
            I => \N__45571\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__45571\,
            I => \N__45567\
        );

    \I__10285\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45564\
        );

    \I__10284\ : Span4Mux_v
    port map (
            O => \N__45567\,
            I => \N__45560\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__45564\,
            I => \N__45557\
        );

    \I__10282\ : InMux
    port map (
            O => \N__45563\,
            I => \N__45554\
        );

    \I__10281\ : Odrv4
    port map (
            O => \N__45560\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__10280\ : Odrv4
    port map (
            O => \N__45557\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__10279\ : LocalMux
    port map (
            O => \N__45554\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__10278\ : InMux
    port map (
            O => \N__45547\,
            I => \N__45544\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__45544\,
            I => \N__45541\
        );

    \I__10276\ : Span4Mux_h
    port map (
            O => \N__45541\,
            I => \N__45538\
        );

    \I__10275\ : Span4Mux_v
    port map (
            O => \N__45538\,
            I => \N__45535\
        );

    \I__10274\ : Odrv4
    port map (
            O => \N__45535\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__10273\ : InMux
    port map (
            O => \N__45532\,
            I => \N__45529\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__45529\,
            I => \N__45526\
        );

    \I__10271\ : Span4Mux_h
    port map (
            O => \N__45526\,
            I => \N__45523\
        );

    \I__10270\ : Span4Mux_v
    port map (
            O => \N__45523\,
            I => \N__45520\
        );

    \I__10269\ : Odrv4
    port map (
            O => \N__45520\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\
        );

    \I__10268\ : InMux
    port map (
            O => \N__45517\,
            I => \N__45513\
        );

    \I__10267\ : InMux
    port map (
            O => \N__45516\,
            I => \N__45510\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__45513\,
            I => \N__45507\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__45510\,
            I => \N__45504\
        );

    \I__10264\ : Span4Mux_v
    port map (
            O => \N__45507\,
            I => \N__45500\
        );

    \I__10263\ : Span4Mux_h
    port map (
            O => \N__45504\,
            I => \N__45497\
        );

    \I__10262\ : InMux
    port map (
            O => \N__45503\,
            I => \N__45494\
        );

    \I__10261\ : Odrv4
    port map (
            O => \N__45500\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10260\ : Odrv4
    port map (
            O => \N__45497\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__45494\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10258\ : CascadeMux
    port map (
            O => \N__45487\,
            I => \N__45484\
        );

    \I__10257\ : InMux
    port map (
            O => \N__45484\,
            I => \N__45481\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__45481\,
            I => \N__45478\
        );

    \I__10255\ : Span4Mux_v
    port map (
            O => \N__45478\,
            I => \N__45475\
        );

    \I__10254\ : Span4Mux_h
    port map (
            O => \N__45475\,
            I => \N__45472\
        );

    \I__10253\ : Odrv4
    port map (
            O => \N__45472\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\
        );

    \I__10252\ : InMux
    port map (
            O => \N__45469\,
            I => \N__45466\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__45466\,
            I => \N__45463\
        );

    \I__10250\ : Span4Mux_h
    port map (
            O => \N__45463\,
            I => \N__45460\
        );

    \I__10249\ : Odrv4
    port map (
            O => \N__45460\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__10248\ : InMux
    port map (
            O => \N__45457\,
            I => \N__45454\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__45454\,
            I => \N__45451\
        );

    \I__10246\ : Span4Mux_v
    port map (
            O => \N__45451\,
            I => \N__45448\
        );

    \I__10245\ : Span4Mux_h
    port map (
            O => \N__45448\,
            I => \N__45445\
        );

    \I__10244\ : Odrv4
    port map (
            O => \N__45445\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__10243\ : InMux
    port map (
            O => \N__45442\,
            I => \N__45437\
        );

    \I__10242\ : InMux
    port map (
            O => \N__45441\,
            I => \N__45434\
        );

    \I__10241\ : InMux
    port map (
            O => \N__45440\,
            I => \N__45431\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__45437\,
            I => \N__45428\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__45434\,
            I => \N__45425\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__45431\,
            I => \N__45422\
        );

    \I__10237\ : Span4Mux_h
    port map (
            O => \N__45428\,
            I => \N__45419\
        );

    \I__10236\ : Span4Mux_v
    port map (
            O => \N__45425\,
            I => \N__45414\
        );

    \I__10235\ : Span4Mux_h
    port map (
            O => \N__45422\,
            I => \N__45414\
        );

    \I__10234\ : Odrv4
    port map (
            O => \N__45419\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__10233\ : Odrv4
    port map (
            O => \N__45414\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__10232\ : InMux
    port map (
            O => \N__45409\,
            I => \N__45406\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__45406\,
            I => \N__45403\
        );

    \I__10230\ : Span4Mux_h
    port map (
            O => \N__45403\,
            I => \N__45400\
        );

    \I__10229\ : Odrv4
    port map (
            O => \N__45400\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__10228\ : InMux
    port map (
            O => \N__45397\,
            I => \N__45394\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__45394\,
            I => \N__45391\
        );

    \I__10226\ : Span4Mux_h
    port map (
            O => \N__45391\,
            I => \N__45387\
        );

    \I__10225\ : CascadeMux
    port map (
            O => \N__45390\,
            I => \N__45383\
        );

    \I__10224\ : Span4Mux_h
    port map (
            O => \N__45387\,
            I => \N__45380\
        );

    \I__10223\ : InMux
    port map (
            O => \N__45386\,
            I => \N__45377\
        );

    \I__10222\ : InMux
    port map (
            O => \N__45383\,
            I => \N__45374\
        );

    \I__10221\ : Odrv4
    port map (
            O => \N__45380\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__45377\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__45374\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10218\ : CascadeMux
    port map (
            O => \N__45367\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__10217\ : InMux
    port map (
            O => \N__45364\,
            I => \N__45361\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__45361\,
            I => \N__45357\
        );

    \I__10215\ : InMux
    port map (
            O => \N__45360\,
            I => \N__45354\
        );

    \I__10214\ : Span4Mux_v
    port map (
            O => \N__45357\,
            I => \N__45351\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__45354\,
            I => \N__45348\
        );

    \I__10212\ : Span4Mux_h
    port map (
            O => \N__45351\,
            I => \N__45343\
        );

    \I__10211\ : Span4Mux_v
    port map (
            O => \N__45348\,
            I => \N__45343\
        );

    \I__10210\ : Odrv4
    port map (
            O => \N__45343\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__10209\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45335\
        );

    \I__10208\ : InMux
    port map (
            O => \N__45339\,
            I => \N__45332\
        );

    \I__10207\ : InMux
    port map (
            O => \N__45338\,
            I => \N__45329\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__45335\,
            I => \N__45324\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__45332\,
            I => \N__45324\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__45329\,
            I => \N__45316\
        );

    \I__10203\ : Span4Mux_h
    port map (
            O => \N__45324\,
            I => \N__45316\
        );

    \I__10202\ : InMux
    port map (
            O => \N__45323\,
            I => \N__45311\
        );

    \I__10201\ : InMux
    port map (
            O => \N__45322\,
            I => \N__45311\
        );

    \I__10200\ : CascadeMux
    port map (
            O => \N__45321\,
            I => \N__45298\
        );

    \I__10199\ : Span4Mux_v
    port map (
            O => \N__45316\,
            I => \N__45291\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__45311\,
            I => \N__45291\
        );

    \I__10197\ : InMux
    port map (
            O => \N__45310\,
            I => \N__45282\
        );

    \I__10196\ : InMux
    port map (
            O => \N__45309\,
            I => \N__45282\
        );

    \I__10195\ : InMux
    port map (
            O => \N__45308\,
            I => \N__45282\
        );

    \I__10194\ : InMux
    port map (
            O => \N__45307\,
            I => \N__45282\
        );

    \I__10193\ : InMux
    port map (
            O => \N__45306\,
            I => \N__45272\
        );

    \I__10192\ : InMux
    port map (
            O => \N__45305\,
            I => \N__45272\
        );

    \I__10191\ : InMux
    port map (
            O => \N__45304\,
            I => \N__45272\
        );

    \I__10190\ : InMux
    port map (
            O => \N__45303\,
            I => \N__45265\
        );

    \I__10189\ : InMux
    port map (
            O => \N__45302\,
            I => \N__45265\
        );

    \I__10188\ : InMux
    port map (
            O => \N__45301\,
            I => \N__45265\
        );

    \I__10187\ : InMux
    port map (
            O => \N__45298\,
            I => \N__45262\
        );

    \I__10186\ : InMux
    port map (
            O => \N__45297\,
            I => \N__45257\
        );

    \I__10185\ : InMux
    port map (
            O => \N__45296\,
            I => \N__45257\
        );

    \I__10184\ : Span4Mux_h
    port map (
            O => \N__45291\,
            I => \N__45252\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__45282\,
            I => \N__45252\
        );

    \I__10182\ : InMux
    port map (
            O => \N__45281\,
            I => \N__45246\
        );

    \I__10181\ : InMux
    port map (
            O => \N__45280\,
            I => \N__45243\
        );

    \I__10180\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45240\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__45272\,
            I => \N__45232\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__45265\,
            I => \N__45229\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__45262\,
            I => \N__45224\
        );

    \I__10176\ : LocalMux
    port map (
            O => \N__45257\,
            I => \N__45224\
        );

    \I__10175\ : Span4Mux_v
    port map (
            O => \N__45252\,
            I => \N__45219\
        );

    \I__10174\ : InMux
    port map (
            O => \N__45251\,
            I => \N__45212\
        );

    \I__10173\ : InMux
    port map (
            O => \N__45250\,
            I => \N__45212\
        );

    \I__10172\ : InMux
    port map (
            O => \N__45249\,
            I => \N__45212\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__45246\,
            I => \N__45208\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__45243\,
            I => \N__45205\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__45240\,
            I => \N__45202\
        );

    \I__10168\ : InMux
    port map (
            O => \N__45239\,
            I => \N__45191\
        );

    \I__10167\ : InMux
    port map (
            O => \N__45238\,
            I => \N__45191\
        );

    \I__10166\ : InMux
    port map (
            O => \N__45237\,
            I => \N__45191\
        );

    \I__10165\ : InMux
    port map (
            O => \N__45236\,
            I => \N__45191\
        );

    \I__10164\ : InMux
    port map (
            O => \N__45235\,
            I => \N__45191\
        );

    \I__10163\ : Span4Mux_h
    port map (
            O => \N__45232\,
            I => \N__45188\
        );

    \I__10162\ : Span4Mux_v
    port map (
            O => \N__45229\,
            I => \N__45183\
        );

    \I__10161\ : Span4Mux_h
    port map (
            O => \N__45224\,
            I => \N__45183\
        );

    \I__10160\ : InMux
    port map (
            O => \N__45223\,
            I => \N__45178\
        );

    \I__10159\ : InMux
    port map (
            O => \N__45222\,
            I => \N__45178\
        );

    \I__10158\ : Sp12to4
    port map (
            O => \N__45219\,
            I => \N__45173\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__45212\,
            I => \N__45173\
        );

    \I__10156\ : InMux
    port map (
            O => \N__45211\,
            I => \N__45170\
        );

    \I__10155\ : Span4Mux_h
    port map (
            O => \N__45208\,
            I => \N__45163\
        );

    \I__10154\ : Span4Mux_v
    port map (
            O => \N__45205\,
            I => \N__45163\
        );

    \I__10153\ : Span4Mux_v
    port map (
            O => \N__45202\,
            I => \N__45163\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__45191\,
            I => \N__45158\
        );

    \I__10151\ : Span4Mux_h
    port map (
            O => \N__45188\,
            I => \N__45158\
        );

    \I__10150\ : Span4Mux_h
    port map (
            O => \N__45183\,
            I => \N__45155\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__45178\,
            I => \N__45150\
        );

    \I__10148\ : Span12Mux_h
    port map (
            O => \N__45173\,
            I => \N__45150\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__45170\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__10146\ : Odrv4
    port map (
            O => \N__45163\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__10145\ : Odrv4
    port map (
            O => \N__45158\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__10144\ : Odrv4
    port map (
            O => \N__45155\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__10143\ : Odrv12
    port map (
            O => \N__45150\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__10142\ : CascadeMux
    port map (
            O => \N__45139\,
            I => \N__45127\
        );

    \I__10141\ : InMux
    port map (
            O => \N__45138\,
            I => \N__45113\
        );

    \I__10140\ : InMux
    port map (
            O => \N__45137\,
            I => \N__45105\
        );

    \I__10139\ : InMux
    port map (
            O => \N__45136\,
            I => \N__45105\
        );

    \I__10138\ : InMux
    port map (
            O => \N__45135\,
            I => \N__45105\
        );

    \I__10137\ : InMux
    port map (
            O => \N__45134\,
            I => \N__45102\
        );

    \I__10136\ : InMux
    port map (
            O => \N__45133\,
            I => \N__45099\
        );

    \I__10135\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45092\
        );

    \I__10134\ : InMux
    port map (
            O => \N__45131\,
            I => \N__45092\
        );

    \I__10133\ : InMux
    port map (
            O => \N__45130\,
            I => \N__45092\
        );

    \I__10132\ : InMux
    port map (
            O => \N__45127\,
            I => \N__45085\
        );

    \I__10131\ : InMux
    port map (
            O => \N__45126\,
            I => \N__45085\
        );

    \I__10130\ : InMux
    port map (
            O => \N__45125\,
            I => \N__45085\
        );

    \I__10129\ : InMux
    port map (
            O => \N__45124\,
            I => \N__45082\
        );

    \I__10128\ : InMux
    port map (
            O => \N__45123\,
            I => \N__45077\
        );

    \I__10127\ : InMux
    port map (
            O => \N__45122\,
            I => \N__45077\
        );

    \I__10126\ : InMux
    port map (
            O => \N__45121\,
            I => \N__45068\
        );

    \I__10125\ : InMux
    port map (
            O => \N__45120\,
            I => \N__45068\
        );

    \I__10124\ : InMux
    port map (
            O => \N__45119\,
            I => \N__45068\
        );

    \I__10123\ : InMux
    port map (
            O => \N__45118\,
            I => \N__45068\
        );

    \I__10122\ : InMux
    port map (
            O => \N__45117\,
            I => \N__45057\
        );

    \I__10121\ : InMux
    port map (
            O => \N__45116\,
            I => \N__45054\
        );

    \I__10120\ : LocalMux
    port map (
            O => \N__45113\,
            I => \N__45051\
        );

    \I__10119\ : InMux
    port map (
            O => \N__45112\,
            I => \N__45048\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__45105\,
            I => \N__45043\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__45102\,
            I => \N__45038\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__45099\,
            I => \N__45038\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__45092\,
            I => \N__45033\
        );

    \I__10114\ : LocalMux
    port map (
            O => \N__45085\,
            I => \N__45033\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__45082\,
            I => \N__45030\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__45077\,
            I => \N__45027\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__45068\,
            I => \N__45024\
        );

    \I__10110\ : InMux
    port map (
            O => \N__45067\,
            I => \N__45021\
        );

    \I__10109\ : InMux
    port map (
            O => \N__45066\,
            I => \N__45016\
        );

    \I__10108\ : InMux
    port map (
            O => \N__45065\,
            I => \N__45016\
        );

    \I__10107\ : InMux
    port map (
            O => \N__45064\,
            I => \N__45005\
        );

    \I__10106\ : InMux
    port map (
            O => \N__45063\,
            I => \N__45005\
        );

    \I__10105\ : InMux
    port map (
            O => \N__45062\,
            I => \N__45005\
        );

    \I__10104\ : InMux
    port map (
            O => \N__45061\,
            I => \N__45005\
        );

    \I__10103\ : InMux
    port map (
            O => \N__45060\,
            I => \N__45005\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__45057\,
            I => \N__45000\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__45054\,
            I => \N__45000\
        );

    \I__10100\ : Span4Mux_h
    port map (
            O => \N__45051\,
            I => \N__44995\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__45048\,
            I => \N__44995\
        );

    \I__10098\ : InMux
    port map (
            O => \N__45047\,
            I => \N__44990\
        );

    \I__10097\ : InMux
    port map (
            O => \N__45046\,
            I => \N__44990\
        );

    \I__10096\ : Span4Mux_v
    port map (
            O => \N__45043\,
            I => \N__44983\
        );

    \I__10095\ : Span4Mux_v
    port map (
            O => \N__45038\,
            I => \N__44983\
        );

    \I__10094\ : Span4Mux_v
    port map (
            O => \N__45033\,
            I => \N__44983\
        );

    \I__10093\ : Span4Mux_v
    port map (
            O => \N__45030\,
            I => \N__44976\
        );

    \I__10092\ : Span4Mux_v
    port map (
            O => \N__45027\,
            I => \N__44976\
        );

    \I__10091\ : Span4Mux_v
    port map (
            O => \N__45024\,
            I => \N__44976\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__45021\,
            I => \N__44973\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__45016\,
            I => \N__44966\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__45005\,
            I => \N__44966\
        );

    \I__10087\ : Span4Mux_h
    port map (
            O => \N__45000\,
            I => \N__44966\
        );

    \I__10086\ : Span4Mux_h
    port map (
            O => \N__44995\,
            I => \N__44963\
        );

    \I__10085\ : LocalMux
    port map (
            O => \N__44990\,
            I => \N__44956\
        );

    \I__10084\ : Sp12to4
    port map (
            O => \N__44983\,
            I => \N__44956\
        );

    \I__10083\ : Sp12to4
    port map (
            O => \N__44976\,
            I => \N__44956\
        );

    \I__10082\ : Odrv4
    port map (
            O => \N__44973\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__10081\ : Odrv4
    port map (
            O => \N__44966\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__10080\ : Odrv4
    port map (
            O => \N__44963\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__10079\ : Odrv12
    port map (
            O => \N__44956\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44947\,
            I => \N__44944\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__44944\,
            I => \N__44941\
        );

    \I__10076\ : Span4Mux_h
    port map (
            O => \N__44941\,
            I => \N__44938\
        );

    \I__10075\ : Odrv4
    port map (
            O => \N__44938\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__10074\ : CascadeMux
    port map (
            O => \N__44935\,
            I => \N__44930\
        );

    \I__10073\ : CascadeMux
    port map (
            O => \N__44934\,
            I => \N__44927\
        );

    \I__10072\ : CascadeMux
    port map (
            O => \N__44933\,
            I => \N__44924\
        );

    \I__10071\ : InMux
    port map (
            O => \N__44930\,
            I => \N__44906\
        );

    \I__10070\ : InMux
    port map (
            O => \N__44927\,
            I => \N__44906\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44924\,
            I => \N__44903\
        );

    \I__10068\ : CascadeMux
    port map (
            O => \N__44923\,
            I => \N__44900\
        );

    \I__10067\ : CascadeMux
    port map (
            O => \N__44922\,
            I => \N__44897\
        );

    \I__10066\ : CascadeMux
    port map (
            O => \N__44921\,
            I => \N__44894\
        );

    \I__10065\ : CascadeMux
    port map (
            O => \N__44920\,
            I => \N__44891\
        );

    \I__10064\ : CascadeMux
    port map (
            O => \N__44919\,
            I => \N__44888\
        );

    \I__10063\ : CascadeMux
    port map (
            O => \N__44918\,
            I => \N__44885\
        );

    \I__10062\ : CascadeMux
    port map (
            O => \N__44917\,
            I => \N__44880\
        );

    \I__10061\ : CascadeMux
    port map (
            O => \N__44916\,
            I => \N__44877\
        );

    \I__10060\ : CascadeMux
    port map (
            O => \N__44915\,
            I => \N__44874\
        );

    \I__10059\ : CascadeMux
    port map (
            O => \N__44914\,
            I => \N__44871\
        );

    \I__10058\ : InMux
    port map (
            O => \N__44913\,
            I => \N__44868\
        );

    \I__10057\ : CascadeMux
    port map (
            O => \N__44912\,
            I => \N__44862\
        );

    \I__10056\ : CascadeMux
    port map (
            O => \N__44911\,
            I => \N__44859\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__44906\,
            I => \N__44856\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__44903\,
            I => \N__44853\
        );

    \I__10053\ : InMux
    port map (
            O => \N__44900\,
            I => \N__44849\
        );

    \I__10052\ : InMux
    port map (
            O => \N__44897\,
            I => \N__44842\
        );

    \I__10051\ : InMux
    port map (
            O => \N__44894\,
            I => \N__44842\
        );

    \I__10050\ : InMux
    port map (
            O => \N__44891\,
            I => \N__44842\
        );

    \I__10049\ : InMux
    port map (
            O => \N__44888\,
            I => \N__44837\
        );

    \I__10048\ : InMux
    port map (
            O => \N__44885\,
            I => \N__44837\
        );

    \I__10047\ : CascadeMux
    port map (
            O => \N__44884\,
            I => \N__44834\
        );

    \I__10046\ : CascadeMux
    port map (
            O => \N__44883\,
            I => \N__44829\
        );

    \I__10045\ : InMux
    port map (
            O => \N__44880\,
            I => \N__44826\
        );

    \I__10044\ : InMux
    port map (
            O => \N__44877\,
            I => \N__44823\
        );

    \I__10043\ : InMux
    port map (
            O => \N__44874\,
            I => \N__44818\
        );

    \I__10042\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44818\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__44868\,
            I => \N__44815\
        );

    \I__10040\ : InMux
    port map (
            O => \N__44867\,
            I => \N__44812\
        );

    \I__10039\ : CascadeMux
    port map (
            O => \N__44866\,
            I => \N__44803\
        );

    \I__10038\ : CascadeMux
    port map (
            O => \N__44865\,
            I => \N__44800\
        );

    \I__10037\ : InMux
    port map (
            O => \N__44862\,
            I => \N__44794\
        );

    \I__10036\ : InMux
    port map (
            O => \N__44859\,
            I => \N__44794\
        );

    \I__10035\ : Span4Mux_h
    port map (
            O => \N__44856\,
            I => \N__44789\
        );

    \I__10034\ : Span4Mux_h
    port map (
            O => \N__44853\,
            I => \N__44789\
        );

    \I__10033\ : InMux
    port map (
            O => \N__44852\,
            I => \N__44786\
        );

    \I__10032\ : LocalMux
    port map (
            O => \N__44849\,
            I => \N__44783\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__44842\,
            I => \N__44778\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__44837\,
            I => \N__44778\
        );

    \I__10029\ : InMux
    port map (
            O => \N__44834\,
            I => \N__44775\
        );

    \I__10028\ : CascadeMux
    port map (
            O => \N__44833\,
            I => \N__44772\
        );

    \I__10027\ : CascadeMux
    port map (
            O => \N__44832\,
            I => \N__44769\
        );

    \I__10026\ : InMux
    port map (
            O => \N__44829\,
            I => \N__44765\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__44826\,
            I => \N__44754\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__44823\,
            I => \N__44754\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__44818\,
            I => \N__44754\
        );

    \I__10022\ : Span4Mux_h
    port map (
            O => \N__44815\,
            I => \N__44754\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__44812\,
            I => \N__44754\
        );

    \I__10020\ : CascadeMux
    port map (
            O => \N__44811\,
            I => \N__44751\
        );

    \I__10019\ : CascadeMux
    port map (
            O => \N__44810\,
            I => \N__44748\
        );

    \I__10018\ : CascadeMux
    port map (
            O => \N__44809\,
            I => \N__44745\
        );

    \I__10017\ : CascadeMux
    port map (
            O => \N__44808\,
            I => \N__44742\
        );

    \I__10016\ : CascadeMux
    port map (
            O => \N__44807\,
            I => \N__44739\
        );

    \I__10015\ : CascadeMux
    port map (
            O => \N__44806\,
            I => \N__44736\
        );

    \I__10014\ : InMux
    port map (
            O => \N__44803\,
            I => \N__44731\
        );

    \I__10013\ : InMux
    port map (
            O => \N__44800\,
            I => \N__44731\
        );

    \I__10012\ : InMux
    port map (
            O => \N__44799\,
            I => \N__44728\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__44794\,
            I => \N__44721\
        );

    \I__10010\ : Span4Mux_v
    port map (
            O => \N__44789\,
            I => \N__44721\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__44786\,
            I => \N__44721\
        );

    \I__10008\ : Span4Mux_v
    port map (
            O => \N__44783\,
            I => \N__44714\
        );

    \I__10007\ : Span4Mux_v
    port map (
            O => \N__44778\,
            I => \N__44714\
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__44775\,
            I => \N__44714\
        );

    \I__10005\ : InMux
    port map (
            O => \N__44772\,
            I => \N__44711\
        );

    \I__10004\ : InMux
    port map (
            O => \N__44769\,
            I => \N__44708\
        );

    \I__10003\ : InMux
    port map (
            O => \N__44768\,
            I => \N__44705\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__44765\,
            I => \N__44702\
        );

    \I__10001\ : Span4Mux_h
    port map (
            O => \N__44754\,
            I => \N__44699\
        );

    \I__10000\ : InMux
    port map (
            O => \N__44751\,
            I => \N__44694\
        );

    \I__9999\ : InMux
    port map (
            O => \N__44748\,
            I => \N__44694\
        );

    \I__9998\ : InMux
    port map (
            O => \N__44745\,
            I => \N__44689\
        );

    \I__9997\ : InMux
    port map (
            O => \N__44742\,
            I => \N__44689\
        );

    \I__9996\ : InMux
    port map (
            O => \N__44739\,
            I => \N__44684\
        );

    \I__9995\ : InMux
    port map (
            O => \N__44736\,
            I => \N__44684\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__44731\,
            I => \N__44675\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__44728\,
            I => \N__44675\
        );

    \I__9992\ : Span4Mux_v
    port map (
            O => \N__44721\,
            I => \N__44675\
        );

    \I__9991\ : Span4Mux_h
    port map (
            O => \N__44714\,
            I => \N__44675\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__44711\,
            I => \N__44664\
        );

    \I__9989\ : LocalMux
    port map (
            O => \N__44708\,
            I => \N__44664\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__44705\,
            I => \N__44664\
        );

    \I__9987\ : Span4Mux_h
    port map (
            O => \N__44702\,
            I => \N__44664\
        );

    \I__9986\ : Span4Mux_h
    port map (
            O => \N__44699\,
            I => \N__44664\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__44694\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__44689\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__44684\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9982\ : Odrv4
    port map (
            O => \N__44675\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9981\ : Odrv4
    port map (
            O => \N__44664\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9980\ : InMux
    port map (
            O => \N__44653\,
            I => \N__44647\
        );

    \I__9979\ : InMux
    port map (
            O => \N__44652\,
            I => \N__44644\
        );

    \I__9978\ : CascadeMux
    port map (
            O => \N__44651\,
            I => \N__44641\
        );

    \I__9977\ : InMux
    port map (
            O => \N__44650\,
            I => \N__44638\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__44647\,
            I => \N__44635\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__44644\,
            I => \N__44632\
        );

    \I__9974\ : InMux
    port map (
            O => \N__44641\,
            I => \N__44629\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__44638\,
            I => \N__44626\
        );

    \I__9972\ : Span4Mux_h
    port map (
            O => \N__44635\,
            I => \N__44622\
        );

    \I__9971\ : Span4Mux_h
    port map (
            O => \N__44632\,
            I => \N__44619\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__44629\,
            I => \N__44614\
        );

    \I__9969\ : Span4Mux_h
    port map (
            O => \N__44626\,
            I => \N__44614\
        );

    \I__9968\ : InMux
    port map (
            O => \N__44625\,
            I => \N__44611\
        );

    \I__9967\ : Span4Mux_h
    port map (
            O => \N__44622\,
            I => \N__44606\
        );

    \I__9966\ : Span4Mux_h
    port map (
            O => \N__44619\,
            I => \N__44606\
        );

    \I__9965\ : Span4Mux_h
    port map (
            O => \N__44614\,
            I => \N__44603\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__44611\,
            I => \N__44600\
        );

    \I__9963\ : Odrv4
    port map (
            O => \N__44606\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__9962\ : Odrv4
    port map (
            O => \N__44603\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__9961\ : Odrv4
    port map (
            O => \N__44600\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__9960\ : CascadeMux
    port map (
            O => \N__44593\,
            I => \N__44590\
        );

    \I__9959\ : InMux
    port map (
            O => \N__44590\,
            I => \N__44587\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__44587\,
            I => \N__44584\
        );

    \I__9957\ : Odrv4
    port map (
            O => \N__44584\,
            I => \current_shift_inst.PI_CTRL.integrator_i_26\
        );

    \I__9956\ : CascadeMux
    port map (
            O => \N__44581\,
            I => \N__44578\
        );

    \I__9955\ : InMux
    port map (
            O => \N__44578\,
            I => \N__44574\
        );

    \I__9954\ : InMux
    port map (
            O => \N__44577\,
            I => \N__44570\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__44574\,
            I => \N__44567\
        );

    \I__9952\ : InMux
    port map (
            O => \N__44573\,
            I => \N__44564\
        );

    \I__9951\ : LocalMux
    port map (
            O => \N__44570\,
            I => \N__44559\
        );

    \I__9950\ : Span4Mux_h
    port map (
            O => \N__44567\,
            I => \N__44556\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__44564\,
            I => \N__44553\
        );

    \I__9948\ : InMux
    port map (
            O => \N__44563\,
            I => \N__44550\
        );

    \I__9947\ : InMux
    port map (
            O => \N__44562\,
            I => \N__44547\
        );

    \I__9946\ : Span4Mux_h
    port map (
            O => \N__44559\,
            I => \N__44544\
        );

    \I__9945\ : Odrv4
    port map (
            O => \N__44556\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__9944\ : Odrv4
    port map (
            O => \N__44553\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__44550\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__9942\ : LocalMux
    port map (
            O => \N__44547\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__9941\ : Odrv4
    port map (
            O => \N__44544\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__9940\ : CascadeMux
    port map (
            O => \N__44533\,
            I => \N__44530\
        );

    \I__9939\ : InMux
    port map (
            O => \N__44530\,
            I => \N__44527\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__44527\,
            I => \N__44524\
        );

    \I__9937\ : Odrv4
    port map (
            O => \N__44524\,
            I => \current_shift_inst.PI_CTRL.integrator_i_24\
        );

    \I__9936\ : InMux
    port map (
            O => \N__44521\,
            I => \N__44517\
        );

    \I__9935\ : CascadeMux
    port map (
            O => \N__44520\,
            I => \N__44514\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__44517\,
            I => \N__44510\
        );

    \I__9933\ : InMux
    port map (
            O => \N__44514\,
            I => \N__44507\
        );

    \I__9932\ : InMux
    port map (
            O => \N__44513\,
            I => \N__44504\
        );

    \I__9931\ : Span4Mux_v
    port map (
            O => \N__44510\,
            I => \N__44501\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__44507\,
            I => \N__44498\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__44504\,
            I => \N__44495\
        );

    \I__9928\ : Span4Mux_h
    port map (
            O => \N__44501\,
            I => \N__44490\
        );

    \I__9927\ : Span4Mux_h
    port map (
            O => \N__44498\,
            I => \N__44490\
        );

    \I__9926\ : Span12Mux_h
    port map (
            O => \N__44495\,
            I => \N__44486\
        );

    \I__9925\ : Span4Mux_h
    port map (
            O => \N__44490\,
            I => \N__44483\
        );

    \I__9924\ : InMux
    port map (
            O => \N__44489\,
            I => \N__44480\
        );

    \I__9923\ : Odrv12
    port map (
            O => \N__44486\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__9922\ : Odrv4
    port map (
            O => \N__44483\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__44480\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__9920\ : CascadeMux
    port map (
            O => \N__44473\,
            I => \N__44470\
        );

    \I__9919\ : InMux
    port map (
            O => \N__44470\,
            I => \N__44467\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__44467\,
            I => \N__44464\
        );

    \I__9917\ : Odrv4
    port map (
            O => \N__44464\,
            I => \current_shift_inst.PI_CTRL.integrator_i_28\
        );

    \I__9916\ : CascadeMux
    port map (
            O => \N__44461\,
            I => \N__44458\
        );

    \I__9915\ : InMux
    port map (
            O => \N__44458\,
            I => \N__44455\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__44455\,
            I => \N__44450\
        );

    \I__9913\ : InMux
    port map (
            O => \N__44454\,
            I => \N__44447\
        );

    \I__9912\ : InMux
    port map (
            O => \N__44453\,
            I => \N__44444\
        );

    \I__9911\ : Span4Mux_v
    port map (
            O => \N__44450\,
            I => \N__44438\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__44447\,
            I => \N__44438\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__44444\,
            I => \N__44435\
        );

    \I__9908\ : InMux
    port map (
            O => \N__44443\,
            I => \N__44432\
        );

    \I__9907\ : Span4Mux_h
    port map (
            O => \N__44438\,
            I => \N__44428\
        );

    \I__9906\ : Span4Mux_h
    port map (
            O => \N__44435\,
            I => \N__44425\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__44432\,
            I => \N__44422\
        );

    \I__9904\ : InMux
    port map (
            O => \N__44431\,
            I => \N__44419\
        );

    \I__9903\ : Span4Mux_h
    port map (
            O => \N__44428\,
            I => \N__44416\
        );

    \I__9902\ : Odrv4
    port map (
            O => \N__44425\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__9901\ : Odrv12
    port map (
            O => \N__44422\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__44419\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__9899\ : Odrv4
    port map (
            O => \N__44416\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__9898\ : CascadeMux
    port map (
            O => \N__44407\,
            I => \N__44404\
        );

    \I__9897\ : InMux
    port map (
            O => \N__44404\,
            I => \N__44401\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__44401\,
            I => \N__44398\
        );

    \I__9895\ : Odrv4
    port map (
            O => \N__44398\,
            I => \current_shift_inst.PI_CTRL.integrator_i_23\
        );

    \I__9894\ : InMux
    port map (
            O => \N__44395\,
            I => \N__44392\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__44392\,
            I => \N__44389\
        );

    \I__9892\ : Span4Mux_h
    port map (
            O => \N__44389\,
            I => \N__44386\
        );

    \I__9891\ : Odrv4
    port map (
            O => \N__44386\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9890\ : InMux
    port map (
            O => \N__44383\,
            I => \N__44380\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__44380\,
            I => \N__44377\
        );

    \I__9888\ : Span4Mux_h
    port map (
            O => \N__44377\,
            I => \N__44374\
        );

    \I__9887\ : Odrv4
    port map (
            O => \N__44374\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9886\ : CascadeMux
    port map (
            O => \N__44371\,
            I => \N__44368\
        );

    \I__9885\ : InMux
    port map (
            O => \N__44368\,
            I => \N__44365\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__44365\,
            I => \N__44362\
        );

    \I__9883\ : Span4Mux_h
    port map (
            O => \N__44362\,
            I => \N__44359\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__44359\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__9881\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44353\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__44353\,
            I => \N__44350\
        );

    \I__9879\ : Span4Mux_v
    port map (
            O => \N__44350\,
            I => \N__44347\
        );

    \I__9878\ : Odrv4
    port map (
            O => \N__44347\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9877\ : InMux
    port map (
            O => \N__44344\,
            I => \N__44341\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__44341\,
            I => \N__44338\
        );

    \I__9875\ : Span12Mux_h
    port map (
            O => \N__44338\,
            I => \N__44335\
        );

    \I__9874\ : Odrv12
    port map (
            O => \N__44335\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\
        );

    \I__9873\ : InMux
    port map (
            O => \N__44332\,
            I => \N__44328\
        );

    \I__9872\ : InMux
    port map (
            O => \N__44331\,
            I => \N__44324\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__44328\,
            I => \N__44321\
        );

    \I__9870\ : InMux
    port map (
            O => \N__44327\,
            I => \N__44318\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__44324\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__9868\ : Odrv4
    port map (
            O => \N__44321\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__44318\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__9866\ : InMux
    port map (
            O => \N__44311\,
            I => \N__44307\
        );

    \I__9865\ : InMux
    port map (
            O => \N__44310\,
            I => \N__44304\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__44307\,
            I => \N__44298\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__44304\,
            I => \N__44298\
        );

    \I__9862\ : InMux
    port map (
            O => \N__44303\,
            I => \N__44295\
        );

    \I__9861\ : Span4Mux_h
    port map (
            O => \N__44298\,
            I => \N__44292\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__44295\,
            I => \N__44289\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__44292\,
            I => \N__44286\
        );

    \I__9858\ : Odrv12
    port map (
            O => \N__44289\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__9857\ : Odrv4
    port map (
            O => \N__44286\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__9856\ : CascadeMux
    port map (
            O => \N__44281\,
            I => \N__44278\
        );

    \I__9855\ : InMux
    port map (
            O => \N__44278\,
            I => \N__44275\
        );

    \I__9854\ : LocalMux
    port map (
            O => \N__44275\,
            I => \N__44272\
        );

    \I__9853\ : Span4Mux_v
    port map (
            O => \N__44272\,
            I => \N__44269\
        );

    \I__9852\ : Odrv4
    port map (
            O => \N__44269\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__9851\ : InMux
    port map (
            O => \N__44266\,
            I => \N__44262\
        );

    \I__9850\ : InMux
    port map (
            O => \N__44265\,
            I => \N__44259\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__44262\,
            I => \N__44256\
        );

    \I__9848\ : LocalMux
    port map (
            O => \N__44259\,
            I => \N__44253\
        );

    \I__9847\ : Span4Mux_h
    port map (
            O => \N__44256\,
            I => \N__44249\
        );

    \I__9846\ : Span12Mux_h
    port map (
            O => \N__44253\,
            I => \N__44246\
        );

    \I__9845\ : InMux
    port map (
            O => \N__44252\,
            I => \N__44243\
        );

    \I__9844\ : Odrv4
    port map (
            O => \N__44249\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__9843\ : Odrv12
    port map (
            O => \N__44246\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__44243\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__9841\ : InMux
    port map (
            O => \N__44236\,
            I => \N__44233\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__44233\,
            I => \N__44230\
        );

    \I__9839\ : Odrv12
    port map (
            O => \N__44230\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_17\
        );

    \I__9838\ : InMux
    port map (
            O => \N__44227\,
            I => \N__44224\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__44224\,
            I => \N__44221\
        );

    \I__9836\ : Odrv4
    port map (
            O => \N__44221\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIKOBPZ0Z_17\
        );

    \I__9835\ : CascadeMux
    port map (
            O => \N__44218\,
            I => \N__44215\
        );

    \I__9834\ : InMux
    port map (
            O => \N__44215\,
            I => \N__44212\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__44212\,
            I => \N__44209\
        );

    \I__9832\ : Span4Mux_h
    port map (
            O => \N__44209\,
            I => \N__44206\
        );

    \I__9831\ : Odrv4
    port map (
            O => \N__44206\,
            I => \current_shift_inst.PI_CTRL.integrator_i_10\
        );

    \I__9830\ : CascadeMux
    port map (
            O => \N__44203\,
            I => \N__44198\
        );

    \I__9829\ : InMux
    port map (
            O => \N__44202\,
            I => \N__44195\
        );

    \I__9828\ : InMux
    port map (
            O => \N__44201\,
            I => \N__44192\
        );

    \I__9827\ : InMux
    port map (
            O => \N__44198\,
            I => \N__44189\
        );

    \I__9826\ : LocalMux
    port map (
            O => \N__44195\,
            I => \N__44186\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__44192\,
            I => \N__44183\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__44189\,
            I => \N__44180\
        );

    \I__9823\ : Span4Mux_h
    port map (
            O => \N__44186\,
            I => \N__44173\
        );

    \I__9822\ : Span4Mux_v
    port map (
            O => \N__44183\,
            I => \N__44173\
        );

    \I__9821\ : Span4Mux_h
    port map (
            O => \N__44180\,
            I => \N__44170\
        );

    \I__9820\ : InMux
    port map (
            O => \N__44179\,
            I => \N__44167\
        );

    \I__9819\ : InMux
    port map (
            O => \N__44178\,
            I => \N__44164\
        );

    \I__9818\ : Span4Mux_h
    port map (
            O => \N__44173\,
            I => \N__44161\
        );

    \I__9817\ : Odrv4
    port map (
            O => \N__44170\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__9816\ : LocalMux
    port map (
            O => \N__44167\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__44164\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__9814\ : Odrv4
    port map (
            O => \N__44161\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__9813\ : CascadeMux
    port map (
            O => \N__44152\,
            I => \N__44149\
        );

    \I__9812\ : InMux
    port map (
            O => \N__44149\,
            I => \N__44146\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__44146\,
            I => \N__44143\
        );

    \I__9810\ : Odrv4
    port map (
            O => \N__44143\,
            I => \current_shift_inst.PI_CTRL.integrator_i_7\
        );

    \I__9809\ : CascadeMux
    port map (
            O => \N__44140\,
            I => \N__44136\
        );

    \I__9808\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44132\
        );

    \I__9807\ : InMux
    port map (
            O => \N__44136\,
            I => \N__44127\
        );

    \I__9806\ : InMux
    port map (
            O => \N__44135\,
            I => \N__44127\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__44132\,
            I => \N__44123\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__44127\,
            I => \N__44120\
        );

    \I__9803\ : CascadeMux
    port map (
            O => \N__44126\,
            I => \N__44116\
        );

    \I__9802\ : Span4Mux_h
    port map (
            O => \N__44123\,
            I => \N__44111\
        );

    \I__9801\ : Span4Mux_h
    port map (
            O => \N__44120\,
            I => \N__44111\
        );

    \I__9800\ : InMux
    port map (
            O => \N__44119\,
            I => \N__44108\
        );

    \I__9799\ : InMux
    port map (
            O => \N__44116\,
            I => \N__44105\
        );

    \I__9798\ : Span4Mux_h
    port map (
            O => \N__44111\,
            I => \N__44102\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__44108\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__44105\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__9795\ : Odrv4
    port map (
            O => \N__44102\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__9794\ : CascadeMux
    port map (
            O => \N__44095\,
            I => \N__44092\
        );

    \I__9793\ : InMux
    port map (
            O => \N__44092\,
            I => \N__44089\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__44089\,
            I => \N__44086\
        );

    \I__9791\ : Odrv4
    port map (
            O => \N__44086\,
            I => \current_shift_inst.PI_CTRL.integrator_i_13\
        );

    \I__9790\ : InMux
    port map (
            O => \N__44083\,
            I => \N__44074\
        );

    \I__9789\ : InMux
    port map (
            O => \N__44082\,
            I => \N__44063\
        );

    \I__9788\ : InMux
    port map (
            O => \N__44081\,
            I => \N__44060\
        );

    \I__9787\ : InMux
    port map (
            O => \N__44080\,
            I => \N__44057\
        );

    \I__9786\ : InMux
    port map (
            O => \N__44079\,
            I => \N__44046\
        );

    \I__9785\ : InMux
    port map (
            O => \N__44078\,
            I => \N__44043\
        );

    \I__9784\ : InMux
    port map (
            O => \N__44077\,
            I => \N__44040\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__44074\,
            I => \N__44037\
        );

    \I__9782\ : InMux
    port map (
            O => \N__44073\,
            I => \N__44020\
        );

    \I__9781\ : InMux
    port map (
            O => \N__44072\,
            I => \N__44020\
        );

    \I__9780\ : InMux
    port map (
            O => \N__44071\,
            I => \N__44020\
        );

    \I__9779\ : InMux
    port map (
            O => \N__44070\,
            I => \N__44020\
        );

    \I__9778\ : InMux
    port map (
            O => \N__44069\,
            I => \N__44020\
        );

    \I__9777\ : InMux
    port map (
            O => \N__44068\,
            I => \N__44020\
        );

    \I__9776\ : InMux
    port map (
            O => \N__44067\,
            I => \N__44020\
        );

    \I__9775\ : InMux
    port map (
            O => \N__44066\,
            I => \N__44020\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__44063\,
            I => \N__44010\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__44060\,
            I => \N__44010\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__44057\,
            I => \N__44010\
        );

    \I__9771\ : InMux
    port map (
            O => \N__44056\,
            I => \N__43999\
        );

    \I__9770\ : InMux
    port map (
            O => \N__44055\,
            I => \N__43999\
        );

    \I__9769\ : InMux
    port map (
            O => \N__44054\,
            I => \N__43999\
        );

    \I__9768\ : InMux
    port map (
            O => \N__44053\,
            I => \N__43999\
        );

    \I__9767\ : InMux
    port map (
            O => \N__44052\,
            I => \N__43999\
        );

    \I__9766\ : InMux
    port map (
            O => \N__44051\,
            I => \N__43993\
        );

    \I__9765\ : InMux
    port map (
            O => \N__44050\,
            I => \N__43988\
        );

    \I__9764\ : InMux
    port map (
            O => \N__44049\,
            I => \N__43988\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__44046\,
            I => \N__43977\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__44043\,
            I => \N__43974\
        );

    \I__9761\ : LocalMux
    port map (
            O => \N__44040\,
            I => \N__43967\
        );

    \I__9760\ : Span4Mux_v
    port map (
            O => \N__44037\,
            I => \N__43967\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__44020\,
            I => \N__43967\
        );

    \I__9758\ : InMux
    port map (
            O => \N__44019\,
            I => \N__43962\
        );

    \I__9757\ : InMux
    port map (
            O => \N__44018\,
            I => \N__43962\
        );

    \I__9756\ : InMux
    port map (
            O => \N__44017\,
            I => \N__43959\
        );

    \I__9755\ : Span4Mux_v
    port map (
            O => \N__44010\,
            I => \N__43954\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__43999\,
            I => \N__43954\
        );

    \I__9753\ : InMux
    port map (
            O => \N__43998\,
            I => \N__43949\
        );

    \I__9752\ : InMux
    port map (
            O => \N__43997\,
            I => \N__43949\
        );

    \I__9751\ : InMux
    port map (
            O => \N__43996\,
            I => \N__43946\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__43993\,
            I => \N__43941\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__43988\,
            I => \N__43941\
        );

    \I__9748\ : InMux
    port map (
            O => \N__43987\,
            I => \N__43928\
        );

    \I__9747\ : InMux
    port map (
            O => \N__43986\,
            I => \N__43928\
        );

    \I__9746\ : InMux
    port map (
            O => \N__43985\,
            I => \N__43928\
        );

    \I__9745\ : InMux
    port map (
            O => \N__43984\,
            I => \N__43928\
        );

    \I__9744\ : InMux
    port map (
            O => \N__43983\,
            I => \N__43928\
        );

    \I__9743\ : InMux
    port map (
            O => \N__43982\,
            I => \N__43928\
        );

    \I__9742\ : InMux
    port map (
            O => \N__43981\,
            I => \N__43923\
        );

    \I__9741\ : InMux
    port map (
            O => \N__43980\,
            I => \N__43923\
        );

    \I__9740\ : Span4Mux_h
    port map (
            O => \N__43977\,
            I => \N__43920\
        );

    \I__9739\ : Span4Mux_v
    port map (
            O => \N__43974\,
            I => \N__43913\
        );

    \I__9738\ : Span4Mux_h
    port map (
            O => \N__43967\,
            I => \N__43913\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__43962\,
            I => \N__43913\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__43959\,
            I => \N__43908\
        );

    \I__9735\ : Span4Mux_h
    port map (
            O => \N__43954\,
            I => \N__43908\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__43949\,
            I => \N__43901\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__43946\,
            I => \N__43901\
        );

    \I__9732\ : Span4Mux_v
    port map (
            O => \N__43941\,
            I => \N__43901\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__43928\,
            I => \N__43898\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__43923\,
            I => \N__43891\
        );

    \I__9729\ : Span4Mux_v
    port map (
            O => \N__43920\,
            I => \N__43891\
        );

    \I__9728\ : Span4Mux_h
    port map (
            O => \N__43913\,
            I => \N__43891\
        );

    \I__9727\ : Span4Mux_v
    port map (
            O => \N__43908\,
            I => \N__43888\
        );

    \I__9726\ : Span4Mux_v
    port map (
            O => \N__43901\,
            I => \N__43885\
        );

    \I__9725\ : Span4Mux_h
    port map (
            O => \N__43898\,
            I => \N__43882\
        );

    \I__9724\ : Odrv4
    port map (
            O => \N__43891\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__9723\ : Odrv4
    port map (
            O => \N__43888\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__9722\ : Odrv4
    port map (
            O => \N__43885\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__9721\ : Odrv4
    port map (
            O => \N__43882\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__9720\ : InMux
    port map (
            O => \N__43873\,
            I => \N__43869\
        );

    \I__9719\ : InMux
    port map (
            O => \N__43872\,
            I => \N__43866\
        );

    \I__9718\ : LocalMux
    port map (
            O => \N__43869\,
            I => \N__43863\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__43866\,
            I => \N__43860\
        );

    \I__9716\ : Span4Mux_v
    port map (
            O => \N__43863\,
            I => \N__43856\
        );

    \I__9715\ : Span4Mux_h
    port map (
            O => \N__43860\,
            I => \N__43853\
        );

    \I__9714\ : InMux
    port map (
            O => \N__43859\,
            I => \N__43850\
        );

    \I__9713\ : Span4Mux_h
    port map (
            O => \N__43856\,
            I => \N__43845\
        );

    \I__9712\ : Span4Mux_h
    port map (
            O => \N__43853\,
            I => \N__43845\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__43850\,
            I => \N__43842\
        );

    \I__9710\ : Odrv4
    port map (
            O => \N__43845\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__9709\ : Odrv4
    port map (
            O => \N__43842\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__9708\ : InMux
    port map (
            O => \N__43837\,
            I => \N__43834\
        );

    \I__9707\ : LocalMux
    port map (
            O => \N__43834\,
            I => \N__43831\
        );

    \I__9706\ : Span4Mux_h
    port map (
            O => \N__43831\,
            I => \N__43828\
        );

    \I__9705\ : Odrv4
    port map (
            O => \N__43828\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_14\
        );

    \I__9704\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43822\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__43822\,
            I => \N__43819\
        );

    \I__9702\ : Span4Mux_v
    port map (
            O => \N__43819\,
            I => \N__43816\
        );

    \I__9701\ : Odrv4
    port map (
            O => \N__43816\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI898PZ0Z_14\
        );

    \I__9700\ : InMux
    port map (
            O => \N__43813\,
            I => \N__43810\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__43810\,
            I => \N__43807\
        );

    \I__9698\ : Span4Mux_h
    port map (
            O => \N__43807\,
            I => \N__43804\
        );

    \I__9697\ : Odrv4
    port map (
            O => \N__43804\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__9696\ : InMux
    port map (
            O => \N__43801\,
            I => \N__43798\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__43798\,
            I => \N__43794\
        );

    \I__9694\ : InMux
    port map (
            O => \N__43797\,
            I => \N__43790\
        );

    \I__9693\ : Span4Mux_v
    port map (
            O => \N__43794\,
            I => \N__43786\
        );

    \I__9692\ : CascadeMux
    port map (
            O => \N__43793\,
            I => \N__43782\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__43790\,
            I => \N__43779\
        );

    \I__9690\ : InMux
    port map (
            O => \N__43789\,
            I => \N__43776\
        );

    \I__9689\ : Span4Mux_h
    port map (
            O => \N__43786\,
            I => \N__43773\
        );

    \I__9688\ : InMux
    port map (
            O => \N__43785\,
            I => \N__43770\
        );

    \I__9687\ : InMux
    port map (
            O => \N__43782\,
            I => \N__43767\
        );

    \I__9686\ : Span12Mux_s9_v
    port map (
            O => \N__43779\,
            I => \N__43762\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__43776\,
            I => \N__43762\
        );

    \I__9684\ : Span4Mux_h
    port map (
            O => \N__43773\,
            I => \N__43757\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__43770\,
            I => \N__43757\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__43767\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__9681\ : Odrv12
    port map (
            O => \N__43762\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__9680\ : Odrv4
    port map (
            O => \N__43757\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__9679\ : InMux
    port map (
            O => \N__43750\,
            I => \N__43747\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__43747\,
            I => \N__43744\
        );

    \I__9677\ : Span4Mux_h
    port map (
            O => \N__43744\,
            I => \N__43741\
        );

    \I__9676\ : Odrv4
    port map (
            O => \N__43741\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__9675\ : InMux
    port map (
            O => \N__43738\,
            I => \N__43735\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__43735\,
            I => \N__43732\
        );

    \I__9673\ : Span4Mux_v
    port map (
            O => \N__43732\,
            I => \N__43729\
        );

    \I__9672\ : Odrv4
    port map (
            O => \N__43729\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__9671\ : InMux
    port map (
            O => \N__43726\,
            I => \N__43723\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__43723\,
            I => \N__43720\
        );

    \I__9669\ : Odrv12
    port map (
            O => \N__43720\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__9668\ : CascadeMux
    port map (
            O => \N__43717\,
            I => \N__43714\
        );

    \I__9667\ : InMux
    port map (
            O => \N__43714\,
            I => \N__43711\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__43711\,
            I => \N__43708\
        );

    \I__9665\ : Odrv4
    port map (
            O => \N__43708\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__9664\ : InMux
    port map (
            O => \N__43705\,
            I => \N__43702\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__43702\,
            I => \N__43698\
        );

    \I__9662\ : InMux
    port map (
            O => \N__43701\,
            I => \N__43695\
        );

    \I__9661\ : Span4Mux_v
    port map (
            O => \N__43698\,
            I => \N__43689\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__43695\,
            I => \N__43689\
        );

    \I__9659\ : InMux
    port map (
            O => \N__43694\,
            I => \N__43686\
        );

    \I__9658\ : Odrv4
    port map (
            O => \N__43689\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__43686\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9656\ : InMux
    port map (
            O => \N__43681\,
            I => \N__43678\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__43678\,
            I => \N__43675\
        );

    \I__9654\ : Odrv12
    port map (
            O => \N__43675\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__9653\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43669\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__43669\,
            I => \N__43666\
        );

    \I__9651\ : Odrv12
    port map (
            O => \N__43666\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__9650\ : InMux
    port map (
            O => \N__43663\,
            I => \N__43658\
        );

    \I__9649\ : InMux
    port map (
            O => \N__43662\,
            I => \N__43654\
        );

    \I__9648\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43651\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__43658\,
            I => \N__43648\
        );

    \I__9646\ : InMux
    port map (
            O => \N__43657\,
            I => \N__43645\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__43654\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__43651\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__9643\ : Odrv12
    port map (
            O => \N__43648\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__43645\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__9641\ : InMux
    port map (
            O => \N__43636\,
            I => \N__43633\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__43633\,
            I => \N__43629\
        );

    \I__9639\ : InMux
    port map (
            O => \N__43632\,
            I => \N__43626\
        );

    \I__9638\ : Span4Mux_v
    port map (
            O => \N__43629\,
            I => \N__43620\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__43626\,
            I => \N__43620\
        );

    \I__9636\ : InMux
    port map (
            O => \N__43625\,
            I => \N__43617\
        );

    \I__9635\ : Span4Mux_h
    port map (
            O => \N__43620\,
            I => \N__43613\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__43617\,
            I => \N__43609\
        );

    \I__9633\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43606\
        );

    \I__9632\ : Span4Mux_h
    port map (
            O => \N__43613\,
            I => \N__43603\
        );

    \I__9631\ : InMux
    port map (
            O => \N__43612\,
            I => \N__43600\
        );

    \I__9630\ : Odrv4
    port map (
            O => \N__43609\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__43606\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__9628\ : Odrv4
    port map (
            O => \N__43603\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__43600\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__9626\ : InMux
    port map (
            O => \N__43591\,
            I => \N__43585\
        );

    \I__9625\ : InMux
    port map (
            O => \N__43590\,
            I => \N__43582\
        );

    \I__9624\ : CascadeMux
    port map (
            O => \N__43589\,
            I => \N__43579\
        );

    \I__9623\ : CascadeMux
    port map (
            O => \N__43588\,
            I => \N__43576\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__43585\,
            I => \N__43573\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__43582\,
            I => \N__43570\
        );

    \I__9620\ : InMux
    port map (
            O => \N__43579\,
            I => \N__43566\
        );

    \I__9619\ : InMux
    port map (
            O => \N__43576\,
            I => \N__43563\
        );

    \I__9618\ : Span12Mux_v
    port map (
            O => \N__43573\,
            I => \N__43560\
        );

    \I__9617\ : Span4Mux_h
    port map (
            O => \N__43570\,
            I => \N__43557\
        );

    \I__9616\ : InMux
    port map (
            O => \N__43569\,
            I => \N__43554\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__43566\,
            I => \N__43551\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__43563\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__9613\ : Odrv12
    port map (
            O => \N__43560\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__9612\ : Odrv4
    port map (
            O => \N__43557\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__43554\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__9610\ : Odrv4
    port map (
            O => \N__43551\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__9609\ : CascadeMux
    port map (
            O => \N__43540\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\
        );

    \I__9608\ : InMux
    port map (
            O => \N__43537\,
            I => \N__43532\
        );

    \I__9607\ : CascadeMux
    port map (
            O => \N__43536\,
            I => \N__43529\
        );

    \I__9606\ : InMux
    port map (
            O => \N__43535\,
            I => \N__43524\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__43532\,
            I => \N__43521\
        );

    \I__9604\ : InMux
    port map (
            O => \N__43529\,
            I => \N__43516\
        );

    \I__9603\ : InMux
    port map (
            O => \N__43528\,
            I => \N__43516\
        );

    \I__9602\ : InMux
    port map (
            O => \N__43527\,
            I => \N__43513\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__43524\,
            I => \N__43508\
        );

    \I__9600\ : Span12Mux_s7_v
    port map (
            O => \N__43521\,
            I => \N__43508\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__43516\,
            I => \N__43505\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__43513\,
            I => \N__43502\
        );

    \I__9597\ : Odrv12
    port map (
            O => \N__43508\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__9596\ : Odrv4
    port map (
            O => \N__43505\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__9595\ : Odrv4
    port map (
            O => \N__43502\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__9594\ : InMux
    port map (
            O => \N__43495\,
            I => \N__43492\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__43492\,
            I => \N__43489\
        );

    \I__9592\ : Odrv12
    port map (
            O => \N__43489\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\
        );

    \I__9591\ : InMux
    port map (
            O => \N__43486\,
            I => \N__43483\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__43483\,
            I => \N__43480\
        );

    \I__9589\ : Odrv4
    port map (
            O => \N__43480\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__9588\ : CascadeMux
    port map (
            O => \N__43477\,
            I => \N__43474\
        );

    \I__9587\ : InMux
    port map (
            O => \N__43474\,
            I => \N__43471\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__43471\,
            I => \N__43465\
        );

    \I__9585\ : InMux
    port map (
            O => \N__43470\,
            I => \N__43462\
        );

    \I__9584\ : InMux
    port map (
            O => \N__43469\,
            I => \N__43459\
        );

    \I__9583\ : InMux
    port map (
            O => \N__43468\,
            I => \N__43456\
        );

    \I__9582\ : Span4Mux_h
    port map (
            O => \N__43465\,
            I => \N__43453\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__43462\,
            I => \N__43447\
        );

    \I__9580\ : LocalMux
    port map (
            O => \N__43459\,
            I => \N__43447\
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__43456\,
            I => \N__43442\
        );

    \I__9578\ : Sp12to4
    port map (
            O => \N__43453\,
            I => \N__43442\
        );

    \I__9577\ : InMux
    port map (
            O => \N__43452\,
            I => \N__43439\
        );

    \I__9576\ : Span12Mux_h
    port map (
            O => \N__43447\,
            I => \N__43436\
        );

    \I__9575\ : Odrv12
    port map (
            O => \N__43442\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__43439\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__9573\ : Odrv12
    port map (
            O => \N__43436\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__9572\ : InMux
    port map (
            O => \N__43429\,
            I => \N__43426\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__43426\,
            I => \N__43423\
        );

    \I__9570\ : Span4Mux_v
    port map (
            O => \N__43423\,
            I => \N__43420\
        );

    \I__9569\ : Odrv4
    port map (
            O => \N__43420\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__9568\ : InMux
    port map (
            O => \N__43417\,
            I => \N__43414\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__43414\,
            I => \N__43411\
        );

    \I__9566\ : Odrv4
    port map (
            O => \N__43411\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__9565\ : InMux
    port map (
            O => \N__43408\,
            I => \N__43405\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__43405\,
            I => \N__43402\
        );

    \I__9563\ : Odrv4
    port map (
            O => \N__43402\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__9562\ : InMux
    port map (
            O => \N__43399\,
            I => \N__43396\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__43396\,
            I => \N__43393\
        );

    \I__9560\ : Odrv4
    port map (
            O => \N__43393\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__9559\ : InMux
    port map (
            O => \N__43390\,
            I => \N__43387\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__43387\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__9557\ : InMux
    port map (
            O => \N__43384\,
            I => \N__43381\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__43381\,
            I => \N__43378\
        );

    \I__9555\ : Odrv4
    port map (
            O => \N__43378\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__9554\ : InMux
    port map (
            O => \N__43375\,
            I => \N__43372\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__43372\,
            I => \N__43368\
        );

    \I__9552\ : InMux
    port map (
            O => \N__43371\,
            I => \N__43365\
        );

    \I__9551\ : Span4Mux_v
    port map (
            O => \N__43368\,
            I => \N__43359\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__43365\,
            I => \N__43359\
        );

    \I__9549\ : InMux
    port map (
            O => \N__43364\,
            I => \N__43356\
        );

    \I__9548\ : Odrv4
    port map (
            O => \N__43359\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__43356\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9546\ : InMux
    port map (
            O => \N__43351\,
            I => \N__43348\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__43348\,
            I => \N__43345\
        );

    \I__9544\ : Odrv12
    port map (
            O => \N__43345\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\
        );

    \I__9543\ : InMux
    port map (
            O => \N__43342\,
            I => \N__43339\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__43339\,
            I => \N__43336\
        );

    \I__9541\ : Odrv4
    port map (
            O => \N__43336\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__9540\ : InMux
    port map (
            O => \N__43333\,
            I => \N__43330\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__43330\,
            I => \N__43327\
        );

    \I__9538\ : Odrv4
    port map (
            O => \N__43327\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__9537\ : InMux
    port map (
            O => \N__43324\,
            I => \N__43321\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__43321\,
            I => \N__43317\
        );

    \I__9535\ : InMux
    port map (
            O => \N__43320\,
            I => \N__43314\
        );

    \I__9534\ : Span4Mux_v
    port map (
            O => \N__43317\,
            I => \N__43308\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__43314\,
            I => \N__43308\
        );

    \I__9532\ : InMux
    port map (
            O => \N__43313\,
            I => \N__43305\
        );

    \I__9531\ : Odrv4
    port map (
            O => \N__43308\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__43305\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9529\ : InMux
    port map (
            O => \N__43300\,
            I => \N__43297\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__43297\,
            I => \N__43294\
        );

    \I__9527\ : Odrv12
    port map (
            O => \N__43294\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__9526\ : InMux
    port map (
            O => \N__43291\,
            I => \bfn_17_18_0_\
        );

    \I__9525\ : InMux
    port map (
            O => \N__43288\,
            I => \N__43284\
        );

    \I__9524\ : InMux
    port map (
            O => \N__43287\,
            I => \N__43281\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__43284\,
            I => \N__43277\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__43281\,
            I => \N__43274\
        );

    \I__9521\ : InMux
    port map (
            O => \N__43280\,
            I => \N__43271\
        );

    \I__9520\ : Span4Mux_h
    port map (
            O => \N__43277\,
            I => \N__43268\
        );

    \I__9519\ : Span4Mux_v
    port map (
            O => \N__43274\,
            I => \N__43263\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__43271\,
            I => \N__43263\
        );

    \I__9517\ : Odrv4
    port map (
            O => \N__43268\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9516\ : Odrv4
    port map (
            O => \N__43263\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9515\ : InMux
    port map (
            O => \N__43258\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__9514\ : InMux
    port map (
            O => \N__43255\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__9513\ : InMux
    port map (
            O => \N__43252\,
            I => \N__43249\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__43249\,
            I => \N__43246\
        );

    \I__9511\ : Span4Mux_v
    port map (
            O => \N__43246\,
            I => \N__43243\
        );

    \I__9510\ : Span4Mux_h
    port map (
            O => \N__43243\,
            I => \N__43238\
        );

    \I__9509\ : InMux
    port map (
            O => \N__43242\,
            I => \N__43233\
        );

    \I__9508\ : InMux
    port map (
            O => \N__43241\,
            I => \N__43233\
        );

    \I__9507\ : Odrv4
    port map (
            O => \N__43238\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__43233\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9505\ : InMux
    port map (
            O => \N__43228\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__9504\ : InMux
    port map (
            O => \N__43225\,
            I => \N__43221\
        );

    \I__9503\ : InMux
    port map (
            O => \N__43224\,
            I => \N__43218\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__43221\,
            I => \N__43212\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__43218\,
            I => \N__43212\
        );

    \I__9500\ : InMux
    port map (
            O => \N__43217\,
            I => \N__43209\
        );

    \I__9499\ : Odrv4
    port map (
            O => \N__43212\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__43209\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9497\ : InMux
    port map (
            O => \N__43204\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__9496\ : InMux
    port map (
            O => \N__43201\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__9495\ : InMux
    port map (
            O => \N__43198\,
            I => \N__43195\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__43195\,
            I => \N__43192\
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__43192\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__9492\ : CascadeMux
    port map (
            O => \N__43189\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\
        );

    \I__9491\ : InMux
    port map (
            O => \N__43186\,
            I => \N__43183\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__43183\,
            I => \N__43180\
        );

    \I__9489\ : Odrv4
    port map (
            O => \N__43180\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__9488\ : InMux
    port map (
            O => \N__43177\,
            I => \N__43174\
        );

    \I__9487\ : LocalMux
    port map (
            O => \N__43174\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__9486\ : InMux
    port map (
            O => \N__43171\,
            I => \N__43167\
        );

    \I__9485\ : InMux
    port map (
            O => \N__43170\,
            I => \N__43164\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__43167\,
            I => \N__43158\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__43164\,
            I => \N__43158\
        );

    \I__9482\ : InMux
    port map (
            O => \N__43163\,
            I => \N__43155\
        );

    \I__9481\ : Odrv4
    port map (
            O => \N__43158\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__43155\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9479\ : CascadeMux
    port map (
            O => \N__43150\,
            I => \N__43147\
        );

    \I__9478\ : InMux
    port map (
            O => \N__43147\,
            I => \N__43144\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__43144\,
            I => \N__43141\
        );

    \I__9476\ : Odrv12
    port map (
            O => \N__43141\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__9475\ : InMux
    port map (
            O => \N__43138\,
            I => \bfn_17_17_0_\
        );

    \I__9474\ : InMux
    port map (
            O => \N__43135\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__9473\ : InMux
    port map (
            O => \N__43132\,
            I => \N__43129\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__43129\,
            I => \N__43124\
        );

    \I__9471\ : InMux
    port map (
            O => \N__43128\,
            I => \N__43119\
        );

    \I__9470\ : InMux
    port map (
            O => \N__43127\,
            I => \N__43119\
        );

    \I__9469\ : Odrv4
    port map (
            O => \N__43124\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__43119\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9467\ : InMux
    port map (
            O => \N__43114\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__9466\ : InMux
    port map (
            O => \N__43111\,
            I => \N__43108\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__43108\,
            I => \N__43103\
        );

    \I__9464\ : InMux
    port map (
            O => \N__43107\,
            I => \N__43098\
        );

    \I__9463\ : InMux
    port map (
            O => \N__43106\,
            I => \N__43098\
        );

    \I__9462\ : Odrv4
    port map (
            O => \N__43103\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__43098\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9460\ : InMux
    port map (
            O => \N__43093\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__9459\ : InMux
    port map (
            O => \N__43090\,
            I => \N__43086\
        );

    \I__9458\ : InMux
    port map (
            O => \N__43089\,
            I => \N__43083\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__43086\,
            I => \N__43080\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__43083\,
            I => \N__43077\
        );

    \I__9455\ : Span4Mux_v
    port map (
            O => \N__43080\,
            I => \N__43071\
        );

    \I__9454\ : Span4Mux_h
    port map (
            O => \N__43077\,
            I => \N__43071\
        );

    \I__9453\ : InMux
    port map (
            O => \N__43076\,
            I => \N__43068\
        );

    \I__9452\ : Odrv4
    port map (
            O => \N__43071\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__43068\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9450\ : InMux
    port map (
            O => \N__43063\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__9449\ : InMux
    port map (
            O => \N__43060\,
            I => \N__43057\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__43057\,
            I => \N__43054\
        );

    \I__9447\ : Span4Mux_v
    port map (
            O => \N__43054\,
            I => \N__43050\
        );

    \I__9446\ : InMux
    port map (
            O => \N__43053\,
            I => \N__43047\
        );

    \I__9445\ : Span4Mux_h
    port map (
            O => \N__43050\,
            I => \N__43042\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__43047\,
            I => \N__43042\
        );

    \I__9443\ : Span4Mux_v
    port map (
            O => \N__43042\,
            I => \N__43038\
        );

    \I__9442\ : InMux
    port map (
            O => \N__43041\,
            I => \N__43035\
        );

    \I__9441\ : Odrv4
    port map (
            O => \N__43038\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__43035\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9439\ : InMux
    port map (
            O => \N__43030\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__9438\ : InMux
    port map (
            O => \N__43027\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__9437\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43021\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__43021\,
            I => \N__43018\
        );

    \I__9435\ : Span4Mux_h
    port map (
            O => \N__43018\,
            I => \N__43013\
        );

    \I__9434\ : InMux
    port map (
            O => \N__43017\,
            I => \N__43008\
        );

    \I__9433\ : InMux
    port map (
            O => \N__43016\,
            I => \N__43008\
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__43013\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__43008\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9430\ : InMux
    port map (
            O => \N__43003\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__9429\ : InMux
    port map (
            O => \N__43000\,
            I => \N__42996\
        );

    \I__9428\ : InMux
    port map (
            O => \N__42999\,
            I => \N__42993\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__42996\,
            I => \N__42990\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__42993\,
            I => \N__42987\
        );

    \I__9425\ : Span4Mux_v
    port map (
            O => \N__42990\,
            I => \N__42981\
        );

    \I__9424\ : Span4Mux_h
    port map (
            O => \N__42987\,
            I => \N__42981\
        );

    \I__9423\ : InMux
    port map (
            O => \N__42986\,
            I => \N__42978\
        );

    \I__9422\ : Odrv4
    port map (
            O => \N__42981\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__42978\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9420\ : InMux
    port map (
            O => \N__42973\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__9419\ : InMux
    port map (
            O => \N__42970\,
            I => \N__42967\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__42967\,
            I => \N__42964\
        );

    \I__9417\ : Span4Mux_h
    port map (
            O => \N__42964\,
            I => \N__42961\
        );

    \I__9416\ : Span4Mux_h
    port map (
            O => \N__42961\,
            I => \N__42956\
        );

    \I__9415\ : InMux
    port map (
            O => \N__42960\,
            I => \N__42953\
        );

    \I__9414\ : InMux
    port map (
            O => \N__42959\,
            I => \N__42950\
        );

    \I__9413\ : Odrv4
    port map (
            O => \N__42956\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__42953\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__42950\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__9410\ : InMux
    port map (
            O => \N__42943\,
            I => \bfn_17_16_0_\
        );

    \I__9409\ : InMux
    port map (
            O => \N__42940\,
            I => \N__42937\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__42937\,
            I => \N__42933\
        );

    \I__9407\ : InMux
    port map (
            O => \N__42936\,
            I => \N__42930\
        );

    \I__9406\ : Span4Mux_v
    port map (
            O => \N__42933\,
            I => \N__42926\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__42930\,
            I => \N__42923\
        );

    \I__9404\ : InMux
    port map (
            O => \N__42929\,
            I => \N__42920\
        );

    \I__9403\ : Odrv4
    port map (
            O => \N__42926\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__9402\ : Odrv12
    port map (
            O => \N__42923\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__42920\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__9400\ : InMux
    port map (
            O => \N__42913\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__9399\ : InMux
    port map (
            O => \N__42910\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__9398\ : InMux
    port map (
            O => \N__42907\,
            I => \N__42904\
        );

    \I__9397\ : LocalMux
    port map (
            O => \N__42904\,
            I => \N__42901\
        );

    \I__9396\ : Span4Mux_h
    port map (
            O => \N__42901\,
            I => \N__42896\
        );

    \I__9395\ : InMux
    port map (
            O => \N__42900\,
            I => \N__42893\
        );

    \I__9394\ : InMux
    port map (
            O => \N__42899\,
            I => \N__42890\
        );

    \I__9393\ : Odrv4
    port map (
            O => \N__42896\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__42893\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__42890\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9390\ : InMux
    port map (
            O => \N__42883\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__9389\ : InMux
    port map (
            O => \N__42880\,
            I => \N__42877\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__42877\,
            I => \N__42873\
        );

    \I__9387\ : InMux
    port map (
            O => \N__42876\,
            I => \N__42870\
        );

    \I__9386\ : Span4Mux_h
    port map (
            O => \N__42873\,
            I => \N__42866\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__42870\,
            I => \N__42863\
        );

    \I__9384\ : InMux
    port map (
            O => \N__42869\,
            I => \N__42860\
        );

    \I__9383\ : Odrv4
    port map (
            O => \N__42866\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9382\ : Odrv4
    port map (
            O => \N__42863\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__42860\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__9380\ : InMux
    port map (
            O => \N__42853\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__9379\ : InMux
    port map (
            O => \N__42850\,
            I => \N__42847\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__42847\,
            I => \N__42843\
        );

    \I__9377\ : InMux
    port map (
            O => \N__42846\,
            I => \N__42840\
        );

    \I__9376\ : Span4Mux_v
    port map (
            O => \N__42843\,
            I => \N__42836\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__42840\,
            I => \N__42833\
        );

    \I__9374\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42830\
        );

    \I__9373\ : Odrv4
    port map (
            O => \N__42836\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9372\ : Odrv12
    port map (
            O => \N__42833\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__42830\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9370\ : InMux
    port map (
            O => \N__42823\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__9369\ : InMux
    port map (
            O => \N__42820\,
            I => \N__42816\
        );

    \I__9368\ : InMux
    port map (
            O => \N__42819\,
            I => \N__42813\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__42816\,
            I => \N__42810\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__42813\,
            I => \N__42807\
        );

    \I__9365\ : Span4Mux_v
    port map (
            O => \N__42810\,
            I => \N__42801\
        );

    \I__9364\ : Span4Mux_h
    port map (
            O => \N__42807\,
            I => \N__42801\
        );

    \I__9363\ : InMux
    port map (
            O => \N__42806\,
            I => \N__42798\
        );

    \I__9362\ : Odrv4
    port map (
            O => \N__42801\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__42798\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9360\ : InMux
    port map (
            O => \N__42793\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__9359\ : InMux
    port map (
            O => \N__42790\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__9358\ : InMux
    port map (
            O => \N__42787\,
            I => \N__42749\
        );

    \I__9357\ : InMux
    port map (
            O => \N__42786\,
            I => \N__42749\
        );

    \I__9356\ : InMux
    port map (
            O => \N__42785\,
            I => \N__42749\
        );

    \I__9355\ : InMux
    port map (
            O => \N__42784\,
            I => \N__42749\
        );

    \I__9354\ : InMux
    port map (
            O => \N__42783\,
            I => \N__42740\
        );

    \I__9353\ : InMux
    port map (
            O => \N__42782\,
            I => \N__42740\
        );

    \I__9352\ : InMux
    port map (
            O => \N__42781\,
            I => \N__42740\
        );

    \I__9351\ : InMux
    port map (
            O => \N__42780\,
            I => \N__42740\
        );

    \I__9350\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42731\
        );

    \I__9349\ : InMux
    port map (
            O => \N__42778\,
            I => \N__42731\
        );

    \I__9348\ : InMux
    port map (
            O => \N__42777\,
            I => \N__42731\
        );

    \I__9347\ : InMux
    port map (
            O => \N__42776\,
            I => \N__42731\
        );

    \I__9346\ : InMux
    port map (
            O => \N__42775\,
            I => \N__42722\
        );

    \I__9345\ : InMux
    port map (
            O => \N__42774\,
            I => \N__42722\
        );

    \I__9344\ : InMux
    port map (
            O => \N__42773\,
            I => \N__42722\
        );

    \I__9343\ : InMux
    port map (
            O => \N__42772\,
            I => \N__42722\
        );

    \I__9342\ : InMux
    port map (
            O => \N__42771\,
            I => \N__42713\
        );

    \I__9341\ : InMux
    port map (
            O => \N__42770\,
            I => \N__42713\
        );

    \I__9340\ : InMux
    port map (
            O => \N__42769\,
            I => \N__42713\
        );

    \I__9339\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42713\
        );

    \I__9338\ : InMux
    port map (
            O => \N__42767\,
            I => \N__42704\
        );

    \I__9337\ : InMux
    port map (
            O => \N__42766\,
            I => \N__42704\
        );

    \I__9336\ : InMux
    port map (
            O => \N__42765\,
            I => \N__42704\
        );

    \I__9335\ : InMux
    port map (
            O => \N__42764\,
            I => \N__42704\
        );

    \I__9334\ : InMux
    port map (
            O => \N__42763\,
            I => \N__42699\
        );

    \I__9333\ : InMux
    port map (
            O => \N__42762\,
            I => \N__42699\
        );

    \I__9332\ : InMux
    port map (
            O => \N__42761\,
            I => \N__42690\
        );

    \I__9331\ : InMux
    port map (
            O => \N__42760\,
            I => \N__42690\
        );

    \I__9330\ : InMux
    port map (
            O => \N__42759\,
            I => \N__42690\
        );

    \I__9329\ : InMux
    port map (
            O => \N__42758\,
            I => \N__42690\
        );

    \I__9328\ : LocalMux
    port map (
            O => \N__42749\,
            I => \N__42687\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__42740\,
            I => \N__42680\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__42731\,
            I => \N__42680\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__42722\,
            I => \N__42680\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__42713\,
            I => \N__42671\
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__42704\,
            I => \N__42671\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__42699\,
            I => \N__42671\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__42690\,
            I => \N__42671\
        );

    \I__9320\ : Span4Mux_v
    port map (
            O => \N__42687\,
            I => \N__42664\
        );

    \I__9319\ : Span4Mux_v
    port map (
            O => \N__42680\,
            I => \N__42664\
        );

    \I__9318\ : Span4Mux_v
    port map (
            O => \N__42671\,
            I => \N__42664\
        );

    \I__9317\ : Span4Mux_v
    port map (
            O => \N__42664\,
            I => \N__42661\
        );

    \I__9316\ : Odrv4
    port map (
            O => \N__42661\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9315\ : InMux
    port map (
            O => \N__42658\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__9314\ : InMux
    port map (
            O => \N__42655\,
            I => \N__42651\
        );

    \I__9313\ : InMux
    port map (
            O => \N__42654\,
            I => \N__42648\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__42651\,
            I => \N__42645\
        );

    \I__9311\ : LocalMux
    port map (
            O => \N__42648\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__9310\ : Odrv4
    port map (
            O => \N__42645\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__9309\ : CEMux
    port map (
            O => \N__42640\,
            I => \N__42635\
        );

    \I__9308\ : CEMux
    port map (
            O => \N__42639\,
            I => \N__42632\
        );

    \I__9307\ : CEMux
    port map (
            O => \N__42638\,
            I => \N__42629\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__42635\,
            I => \N__42624\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__42632\,
            I => \N__42624\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__42629\,
            I => \N__42620\
        );

    \I__9303\ : Span4Mux_v
    port map (
            O => \N__42624\,
            I => \N__42617\
        );

    \I__9302\ : CEMux
    port map (
            O => \N__42623\,
            I => \N__42614\
        );

    \I__9301\ : Span4Mux_v
    port map (
            O => \N__42620\,
            I => \N__42607\
        );

    \I__9300\ : Span4Mux_h
    port map (
            O => \N__42617\,
            I => \N__42607\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__42614\,
            I => \N__42607\
        );

    \I__9298\ : Span4Mux_v
    port map (
            O => \N__42607\,
            I => \N__42604\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__42604\,
            I => \delay_measurement_inst.delay_tr_timer.N_305_i\
        );

    \I__9296\ : InMux
    port map (
            O => \N__42601\,
            I => \N__42598\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__42598\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__9294\ : CascadeMux
    port map (
            O => \N__42595\,
            I => \N__42592\
        );

    \I__9293\ : InMux
    port map (
            O => \N__42592\,
            I => \N__42583\
        );

    \I__9292\ : InMux
    port map (
            O => \N__42591\,
            I => \N__42583\
        );

    \I__9291\ : InMux
    port map (
            O => \N__42590\,
            I => \N__42583\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__42583\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__9289\ : InMux
    port map (
            O => \N__42580\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__9288\ : InMux
    port map (
            O => \N__42577\,
            I => \N__42568\
        );

    \I__9287\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42568\
        );

    \I__9286\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42568\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__42568\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__9284\ : InMux
    port map (
            O => \N__42565\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__9283\ : InMux
    port map (
            O => \N__42562\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__9282\ : InMux
    port map (
            O => \N__42559\,
            I => \N__42555\
        );

    \I__9281\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42552\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__42555\,
            I => \N__42548\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__42552\,
            I => \N__42545\
        );

    \I__9278\ : InMux
    port map (
            O => \N__42551\,
            I => \N__42542\
        );

    \I__9277\ : Odrv4
    port map (
            O => \N__42548\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__9276\ : Odrv12
    port map (
            O => \N__42545\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__42542\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__9274\ : InMux
    port map (
            O => \N__42535\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__9273\ : InMux
    port map (
            O => \N__42532\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__9272\ : InMux
    port map (
            O => \N__42529\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__9271\ : InMux
    port map (
            O => \N__42526\,
            I => \N__42519\
        );

    \I__9270\ : InMux
    port map (
            O => \N__42525\,
            I => \N__42519\
        );

    \I__9269\ : InMux
    port map (
            O => \N__42524\,
            I => \N__42516\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__42519\,
            I => \N__42513\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__42516\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__9266\ : Odrv4
    port map (
            O => \N__42513\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__9265\ : InMux
    port map (
            O => \N__42508\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__9264\ : InMux
    port map (
            O => \N__42505\,
            I => \N__42498\
        );

    \I__9263\ : InMux
    port map (
            O => \N__42504\,
            I => \N__42498\
        );

    \I__9262\ : InMux
    port map (
            O => \N__42503\,
            I => \N__42495\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__42498\,
            I => \N__42492\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__42495\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__9259\ : Odrv12
    port map (
            O => \N__42492\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__9258\ : InMux
    port map (
            O => \N__42487\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__9257\ : CascadeMux
    port map (
            O => \N__42484\,
            I => \N__42480\
        );

    \I__9256\ : CascadeMux
    port map (
            O => \N__42483\,
            I => \N__42477\
        );

    \I__9255\ : InMux
    port map (
            O => \N__42480\,
            I => \N__42471\
        );

    \I__9254\ : InMux
    port map (
            O => \N__42477\,
            I => \N__42471\
        );

    \I__9253\ : InMux
    port map (
            O => \N__42476\,
            I => \N__42468\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__42471\,
            I => \N__42465\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__42468\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__9250\ : Odrv12
    port map (
            O => \N__42465\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__9249\ : InMux
    port map (
            O => \N__42460\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__9248\ : CascadeMux
    port map (
            O => \N__42457\,
            I => \N__42453\
        );

    \I__9247\ : CascadeMux
    port map (
            O => \N__42456\,
            I => \N__42450\
        );

    \I__9246\ : InMux
    port map (
            O => \N__42453\,
            I => \N__42444\
        );

    \I__9245\ : InMux
    port map (
            O => \N__42450\,
            I => \N__42444\
        );

    \I__9244\ : InMux
    port map (
            O => \N__42449\,
            I => \N__42441\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__42444\,
            I => \N__42438\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__42441\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__9241\ : Odrv12
    port map (
            O => \N__42438\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__9240\ : InMux
    port map (
            O => \N__42433\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__9239\ : InMux
    port map (
            O => \N__42430\,
            I => \N__42426\
        );

    \I__9238\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42422\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__42426\,
            I => \N__42419\
        );

    \I__9236\ : InMux
    port map (
            O => \N__42425\,
            I => \N__42416\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__42422\,
            I => \N__42411\
        );

    \I__9234\ : Span4Mux_v
    port map (
            O => \N__42419\,
            I => \N__42411\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__42416\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__9232\ : Odrv4
    port map (
            O => \N__42411\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__9231\ : InMux
    port map (
            O => \N__42406\,
            I => \bfn_17_14_0_\
        );

    \I__9230\ : InMux
    port map (
            O => \N__42403\,
            I => \N__42399\
        );

    \I__9229\ : InMux
    port map (
            O => \N__42402\,
            I => \N__42396\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__42399\,
            I => \N__42393\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__42396\,
            I => \N__42387\
        );

    \I__9226\ : Span4Mux_v
    port map (
            O => \N__42393\,
            I => \N__42387\
        );

    \I__9225\ : InMux
    port map (
            O => \N__42392\,
            I => \N__42384\
        );

    \I__9224\ : Span4Mux_h
    port map (
            O => \N__42387\,
            I => \N__42381\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__42384\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__9222\ : Odrv4
    port map (
            O => \N__42381\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__9221\ : InMux
    port map (
            O => \N__42376\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__9220\ : CascadeMux
    port map (
            O => \N__42373\,
            I => \N__42369\
        );

    \I__9219\ : CascadeMux
    port map (
            O => \N__42372\,
            I => \N__42366\
        );

    \I__9218\ : InMux
    port map (
            O => \N__42369\,
            I => \N__42360\
        );

    \I__9217\ : InMux
    port map (
            O => \N__42366\,
            I => \N__42360\
        );

    \I__9216\ : InMux
    port map (
            O => \N__42365\,
            I => \N__42357\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__42360\,
            I => \N__42354\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__42357\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__9213\ : Odrv4
    port map (
            O => \N__42354\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__9212\ : InMux
    port map (
            O => \N__42349\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__9211\ : CascadeMux
    port map (
            O => \N__42346\,
            I => \N__42342\
        );

    \I__9210\ : CascadeMux
    port map (
            O => \N__42345\,
            I => \N__42339\
        );

    \I__9209\ : InMux
    port map (
            O => \N__42342\,
            I => \N__42333\
        );

    \I__9208\ : InMux
    port map (
            O => \N__42339\,
            I => \N__42333\
        );

    \I__9207\ : InMux
    port map (
            O => \N__42338\,
            I => \N__42330\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__42333\,
            I => \N__42327\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__42330\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__9204\ : Odrv4
    port map (
            O => \N__42327\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__9203\ : InMux
    port map (
            O => \N__42322\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__9202\ : InMux
    port map (
            O => \N__42319\,
            I => \N__42315\
        );

    \I__9201\ : InMux
    port map (
            O => \N__42318\,
            I => \N__42312\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__42315\,
            I => \N__42309\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__42312\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__9198\ : Odrv12
    port map (
            O => \N__42309\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__9197\ : InMux
    port map (
            O => \N__42304\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__9196\ : InMux
    port map (
            O => \N__42301\,
            I => \N__42295\
        );

    \I__9195\ : InMux
    port map (
            O => \N__42300\,
            I => \N__42295\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__42295\,
            I => \N__42291\
        );

    \I__9193\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42288\
        );

    \I__9192\ : Span4Mux_h
    port map (
            O => \N__42291\,
            I => \N__42285\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__42288\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__9190\ : Odrv4
    port map (
            O => \N__42285\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__9189\ : InMux
    port map (
            O => \N__42280\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__9188\ : InMux
    port map (
            O => \N__42277\,
            I => \N__42270\
        );

    \I__9187\ : InMux
    port map (
            O => \N__42276\,
            I => \N__42270\
        );

    \I__9186\ : InMux
    port map (
            O => \N__42275\,
            I => \N__42267\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__42270\,
            I => \N__42264\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__42267\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__9183\ : Odrv4
    port map (
            O => \N__42264\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__9182\ : InMux
    port map (
            O => \N__42259\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__9181\ : CascadeMux
    port map (
            O => \N__42256\,
            I => \N__42252\
        );

    \I__9180\ : CascadeMux
    port map (
            O => \N__42255\,
            I => \N__42249\
        );

    \I__9179\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42243\
        );

    \I__9178\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42243\
        );

    \I__9177\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42240\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__42243\,
            I => \N__42237\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__42240\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__9174\ : Odrv12
    port map (
            O => \N__42237\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__9173\ : InMux
    port map (
            O => \N__42232\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__9172\ : CascadeMux
    port map (
            O => \N__42229\,
            I => \N__42225\
        );

    \I__9171\ : CascadeMux
    port map (
            O => \N__42228\,
            I => \N__42222\
        );

    \I__9170\ : InMux
    port map (
            O => \N__42225\,
            I => \N__42216\
        );

    \I__9169\ : InMux
    port map (
            O => \N__42222\,
            I => \N__42216\
        );

    \I__9168\ : InMux
    port map (
            O => \N__42221\,
            I => \N__42213\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__42216\,
            I => \N__42210\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__42213\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__9165\ : Odrv12
    port map (
            O => \N__42210\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__9164\ : InMux
    port map (
            O => \N__42205\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__9163\ : InMux
    port map (
            O => \N__42202\,
            I => \N__42198\
        );

    \I__9162\ : InMux
    port map (
            O => \N__42201\,
            I => \N__42195\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__42198\,
            I => \N__42192\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__42195\,
            I => \N__42186\
        );

    \I__9159\ : Span4Mux_v
    port map (
            O => \N__42192\,
            I => \N__42186\
        );

    \I__9158\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42183\
        );

    \I__9157\ : Span4Mux_h
    port map (
            O => \N__42186\,
            I => \N__42180\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__42183\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__9155\ : Odrv4
    port map (
            O => \N__42180\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__9154\ : InMux
    port map (
            O => \N__42175\,
            I => \bfn_17_13_0_\
        );

    \I__9153\ : InMux
    port map (
            O => \N__42172\,
            I => \N__42168\
        );

    \I__9152\ : InMux
    port map (
            O => \N__42171\,
            I => \N__42164\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__42168\,
            I => \N__42161\
        );

    \I__9150\ : InMux
    port map (
            O => \N__42167\,
            I => \N__42158\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__42164\,
            I => \N__42153\
        );

    \I__9148\ : Span4Mux_v
    port map (
            O => \N__42161\,
            I => \N__42153\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__42158\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__9146\ : Odrv4
    port map (
            O => \N__42153\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__9145\ : InMux
    port map (
            O => \N__42148\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__9144\ : CascadeMux
    port map (
            O => \N__42145\,
            I => \N__42141\
        );

    \I__9143\ : CascadeMux
    port map (
            O => \N__42144\,
            I => \N__42138\
        );

    \I__9142\ : InMux
    port map (
            O => \N__42141\,
            I => \N__42132\
        );

    \I__9141\ : InMux
    port map (
            O => \N__42138\,
            I => \N__42132\
        );

    \I__9140\ : InMux
    port map (
            O => \N__42137\,
            I => \N__42129\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__42132\,
            I => \N__42126\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__42129\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__9137\ : Odrv4
    port map (
            O => \N__42126\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__9136\ : InMux
    port map (
            O => \N__42121\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__9135\ : CascadeMux
    port map (
            O => \N__42118\,
            I => \N__42114\
        );

    \I__9134\ : CascadeMux
    port map (
            O => \N__42117\,
            I => \N__42111\
        );

    \I__9133\ : InMux
    port map (
            O => \N__42114\,
            I => \N__42105\
        );

    \I__9132\ : InMux
    port map (
            O => \N__42111\,
            I => \N__42105\
        );

    \I__9131\ : InMux
    port map (
            O => \N__42110\,
            I => \N__42102\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__42105\,
            I => \N__42099\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__42102\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__9128\ : Odrv4
    port map (
            O => \N__42099\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__9127\ : InMux
    port map (
            O => \N__42094\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__9126\ : CascadeMux
    port map (
            O => \N__42091\,
            I => \N__42087\
        );

    \I__9125\ : CascadeMux
    port map (
            O => \N__42090\,
            I => \N__42084\
        );

    \I__9124\ : InMux
    port map (
            O => \N__42087\,
            I => \N__42078\
        );

    \I__9123\ : InMux
    port map (
            O => \N__42084\,
            I => \N__42078\
        );

    \I__9122\ : InMux
    port map (
            O => \N__42083\,
            I => \N__42075\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__42078\,
            I => \N__42072\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__42075\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__9119\ : Odrv12
    port map (
            O => \N__42072\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__9118\ : InMux
    port map (
            O => \N__42067\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__9117\ : InMux
    port map (
            O => \N__42064\,
            I => \N__42057\
        );

    \I__9116\ : InMux
    port map (
            O => \N__42063\,
            I => \N__42057\
        );

    \I__9115\ : InMux
    port map (
            O => \N__42062\,
            I => \N__42054\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__42057\,
            I => \N__42051\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__42054\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__9112\ : Odrv12
    port map (
            O => \N__42051\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__9111\ : InMux
    port map (
            O => \N__42046\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__9110\ : InMux
    port map (
            O => \N__42043\,
            I => \N__42037\
        );

    \I__9109\ : InMux
    port map (
            O => \N__42042\,
            I => \N__42037\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__42037\,
            I => \N__42033\
        );

    \I__9107\ : InMux
    port map (
            O => \N__42036\,
            I => \N__42030\
        );

    \I__9106\ : Span4Mux_h
    port map (
            O => \N__42033\,
            I => \N__42027\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__42030\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__9104\ : Odrv4
    port map (
            O => \N__42027\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__9103\ : InMux
    port map (
            O => \N__42022\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__9102\ : CascadeMux
    port map (
            O => \N__42019\,
            I => \N__42015\
        );

    \I__9101\ : CascadeMux
    port map (
            O => \N__42018\,
            I => \N__42012\
        );

    \I__9100\ : InMux
    port map (
            O => \N__42015\,
            I => \N__42006\
        );

    \I__9099\ : InMux
    port map (
            O => \N__42012\,
            I => \N__42006\
        );

    \I__9098\ : InMux
    port map (
            O => \N__42011\,
            I => \N__42003\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__42006\,
            I => \N__42000\
        );

    \I__9096\ : LocalMux
    port map (
            O => \N__42003\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__9095\ : Odrv12
    port map (
            O => \N__42000\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__9094\ : InMux
    port map (
            O => \N__41995\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__9093\ : CascadeMux
    port map (
            O => \N__41992\,
            I => \N__41988\
        );

    \I__9092\ : CascadeMux
    port map (
            O => \N__41991\,
            I => \N__41985\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41988\,
            I => \N__41979\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41985\,
            I => \N__41979\
        );

    \I__9089\ : InMux
    port map (
            O => \N__41984\,
            I => \N__41976\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__41979\,
            I => \N__41973\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__41976\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__9086\ : Odrv4
    port map (
            O => \N__41973\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__9085\ : InMux
    port map (
            O => \N__41968\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41965\,
            I => \N__41961\
        );

    \I__9083\ : InMux
    port map (
            O => \N__41964\,
            I => \N__41957\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__41961\,
            I => \N__41954\
        );

    \I__9081\ : InMux
    port map (
            O => \N__41960\,
            I => \N__41951\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__41957\,
            I => \N__41946\
        );

    \I__9079\ : Span4Mux_v
    port map (
            O => \N__41954\,
            I => \N__41946\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__41951\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__9077\ : Odrv4
    port map (
            O => \N__41946\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41941\,
            I => \bfn_17_12_0_\
        );

    \I__9075\ : InMux
    port map (
            O => \N__41938\,
            I => \N__41934\
        );

    \I__9074\ : InMux
    port map (
            O => \N__41937\,
            I => \N__41931\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__41934\,
            I => \N__41928\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__41931\,
            I => \N__41922\
        );

    \I__9071\ : Span4Mux_v
    port map (
            O => \N__41928\,
            I => \N__41922\
        );

    \I__9070\ : InMux
    port map (
            O => \N__41927\,
            I => \N__41919\
        );

    \I__9069\ : Span4Mux_h
    port map (
            O => \N__41922\,
            I => \N__41916\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__41919\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__9067\ : Odrv4
    port map (
            O => \N__41916\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__9066\ : InMux
    port map (
            O => \N__41911\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__9065\ : CascadeMux
    port map (
            O => \N__41908\,
            I => \N__41904\
        );

    \I__9064\ : CascadeMux
    port map (
            O => \N__41907\,
            I => \N__41901\
        );

    \I__9063\ : InMux
    port map (
            O => \N__41904\,
            I => \N__41895\
        );

    \I__9062\ : InMux
    port map (
            O => \N__41901\,
            I => \N__41895\
        );

    \I__9061\ : InMux
    port map (
            O => \N__41900\,
            I => \N__41892\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__41895\,
            I => \N__41889\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__41892\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__9058\ : Odrv4
    port map (
            O => \N__41889\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__9057\ : InMux
    port map (
            O => \N__41884\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__9056\ : CascadeMux
    port map (
            O => \N__41881\,
            I => \N__41877\
        );

    \I__9055\ : CascadeMux
    port map (
            O => \N__41880\,
            I => \N__41874\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41877\,
            I => \N__41868\
        );

    \I__9053\ : InMux
    port map (
            O => \N__41874\,
            I => \N__41868\
        );

    \I__9052\ : InMux
    port map (
            O => \N__41873\,
            I => \N__41865\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__41868\,
            I => \N__41862\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__41865\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__9049\ : Odrv4
    port map (
            O => \N__41862\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__9048\ : InMux
    port map (
            O => \N__41857\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__9047\ : InMux
    port map (
            O => \N__41854\,
            I => \N__41851\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__41851\,
            I => \N__41848\
        );

    \I__9045\ : Span4Mux_v
    port map (
            O => \N__41848\,
            I => \N__41845\
        );

    \I__9044\ : Odrv4
    port map (
            O => \N__41845\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_21\
        );

    \I__9043\ : InMux
    port map (
            O => \N__41842\,
            I => \N__41838\
        );

    \I__9042\ : InMux
    port map (
            O => \N__41841\,
            I => \N__41835\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__41838\,
            I => \N__41832\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__41835\,
            I => \N__41829\
        );

    \I__9039\ : Span4Mux_h
    port map (
            O => \N__41832\,
            I => \N__41825\
        );

    \I__9038\ : Span4Mux_h
    port map (
            O => \N__41829\,
            I => \N__41822\
        );

    \I__9037\ : InMux
    port map (
            O => \N__41828\,
            I => \N__41819\
        );

    \I__9036\ : Odrv4
    port map (
            O => \N__41825\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__9035\ : Odrv4
    port map (
            O => \N__41822\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__41819\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__9033\ : InMux
    port map (
            O => \N__41812\,
            I => \N__41809\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__41809\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI9BAQZ0Z_21\
        );

    \I__9031\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41803\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__41803\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__9029\ : CascadeMux
    port map (
            O => \N__41800\,
            I => \N__41796\
        );

    \I__9028\ : InMux
    port map (
            O => \N__41799\,
            I => \N__41793\
        );

    \I__9027\ : InMux
    port map (
            O => \N__41796\,
            I => \N__41790\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__41793\,
            I => \N__41786\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__41790\,
            I => \N__41783\
        );

    \I__9024\ : InMux
    port map (
            O => \N__41789\,
            I => \N__41780\
        );

    \I__9023\ : Span4Mux_v
    port map (
            O => \N__41786\,
            I => \N__41775\
        );

    \I__9022\ : Span4Mux_h
    port map (
            O => \N__41783\,
            I => \N__41770\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__41780\,
            I => \N__41770\
        );

    \I__9020\ : InMux
    port map (
            O => \N__41779\,
            I => \N__41767\
        );

    \I__9019\ : CascadeMux
    port map (
            O => \N__41778\,
            I => \N__41764\
        );

    \I__9018\ : Span4Mux_h
    port map (
            O => \N__41775\,
            I => \N__41757\
        );

    \I__9017\ : Span4Mux_v
    port map (
            O => \N__41770\,
            I => \N__41757\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__41767\,
            I => \N__41757\
        );

    \I__9015\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41754\
        );

    \I__9014\ : Span4Mux_h
    port map (
            O => \N__41757\,
            I => \N__41751\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__41754\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__9012\ : Odrv4
    port map (
            O => \N__41751\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__9011\ : InMux
    port map (
            O => \N__41746\,
            I => \N__41743\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__41743\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__9009\ : CascadeMux
    port map (
            O => \N__41740\,
            I => \N__41736\
        );

    \I__9008\ : InMux
    port map (
            O => \N__41739\,
            I => \N__41733\
        );

    \I__9007\ : InMux
    port map (
            O => \N__41736\,
            I => \N__41730\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__41733\,
            I => \N__41725\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__41730\,
            I => \N__41722\
        );

    \I__9004\ : InMux
    port map (
            O => \N__41729\,
            I => \N__41719\
        );

    \I__9003\ : InMux
    port map (
            O => \N__41728\,
            I => \N__41715\
        );

    \I__9002\ : Span4Mux_v
    port map (
            O => \N__41725\,
            I => \N__41712\
        );

    \I__9001\ : Span4Mux_v
    port map (
            O => \N__41722\,
            I => \N__41709\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__41719\,
            I => \N__41706\
        );

    \I__8999\ : InMux
    port map (
            O => \N__41718\,
            I => \N__41703\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__41715\,
            I => \N__41700\
        );

    \I__8997\ : Span4Mux_h
    port map (
            O => \N__41712\,
            I => \N__41691\
        );

    \I__8996\ : Span4Mux_h
    port map (
            O => \N__41709\,
            I => \N__41691\
        );

    \I__8995\ : Span4Mux_v
    port map (
            O => \N__41706\,
            I => \N__41691\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__41703\,
            I => \N__41691\
        );

    \I__8993\ : Span4Mux_h
    port map (
            O => \N__41700\,
            I => \N__41688\
        );

    \I__8992\ : Span4Mux_h
    port map (
            O => \N__41691\,
            I => \N__41685\
        );

    \I__8991\ : Odrv4
    port map (
            O => \N__41688\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__8990\ : Odrv4
    port map (
            O => \N__41685\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__8989\ : InMux
    port map (
            O => \N__41680\,
            I => \N__41677\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__41677\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__8987\ : CascadeMux
    port map (
            O => \N__41674\,
            I => \N__41671\
        );

    \I__8986\ : InMux
    port map (
            O => \N__41671\,
            I => \N__41667\
        );

    \I__8985\ : InMux
    port map (
            O => \N__41670\,
            I => \N__41664\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__41667\,
            I => \N__41659\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__41664\,
            I => \N__41656\
        );

    \I__8982\ : InMux
    port map (
            O => \N__41663\,
            I => \N__41651\
        );

    \I__8981\ : InMux
    port map (
            O => \N__41662\,
            I => \N__41651\
        );

    \I__8980\ : Span4Mux_h
    port map (
            O => \N__41659\,
            I => \N__41644\
        );

    \I__8979\ : Span4Mux_h
    port map (
            O => \N__41656\,
            I => \N__41644\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__41651\,
            I => \N__41644\
        );

    \I__8977\ : Span4Mux_h
    port map (
            O => \N__41644\,
            I => \N__41641\
        );

    \I__8976\ : Span4Mux_h
    port map (
            O => \N__41641\,
            I => \N__41637\
        );

    \I__8975\ : InMux
    port map (
            O => \N__41640\,
            I => \N__41634\
        );

    \I__8974\ : Odrv4
    port map (
            O => \N__41637\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__41634\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__8972\ : CascadeMux
    port map (
            O => \N__41629\,
            I => \N__41626\
        );

    \I__8971\ : InMux
    port map (
            O => \N__41626\,
            I => \N__41623\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__41623\,
            I => \N__41620\
        );

    \I__8969\ : Odrv4
    port map (
            O => \N__41620\,
            I => \current_shift_inst.PI_CTRL.integrator_i_12\
        );

    \I__8968\ : InMux
    port map (
            O => \N__41617\,
            I => \bfn_17_11_0_\
        );

    \I__8967\ : InMux
    port map (
            O => \N__41614\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__8966\ : CascadeMux
    port map (
            O => \N__41611\,
            I => \N__41607\
        );

    \I__8965\ : CascadeMux
    port map (
            O => \N__41610\,
            I => \N__41604\
        );

    \I__8964\ : InMux
    port map (
            O => \N__41607\,
            I => \N__41598\
        );

    \I__8963\ : InMux
    port map (
            O => \N__41604\,
            I => \N__41598\
        );

    \I__8962\ : InMux
    port map (
            O => \N__41603\,
            I => \N__41595\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__41598\,
            I => \N__41592\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__41595\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8959\ : Odrv4
    port map (
            O => \N__41592\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8958\ : InMux
    port map (
            O => \N__41587\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__8957\ : InMux
    port map (
            O => \N__41584\,
            I => \N__41581\
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__41581\,
            I => \N__41578\
        );

    \I__8955\ : Span4Mux_h
    port map (
            O => \N__41578\,
            I => \N__41575\
        );

    \I__8954\ : Odrv4
    port map (
            O => \N__41575\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__8953\ : InMux
    port map (
            O => \N__41572\,
            I => \N__41568\
        );

    \I__8952\ : InMux
    port map (
            O => \N__41571\,
            I => \N__41565\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__41568\,
            I => \N__41562\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__41565\,
            I => \N__41559\
        );

    \I__8949\ : Span4Mux_h
    port map (
            O => \N__41562\,
            I => \N__41555\
        );

    \I__8948\ : Span4Mux_h
    port map (
            O => \N__41559\,
            I => \N__41552\
        );

    \I__8947\ : InMux
    port map (
            O => \N__41558\,
            I => \N__41549\
        );

    \I__8946\ : Odrv4
    port map (
            O => \N__41555\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__8945\ : Odrv4
    port map (
            O => \N__41552\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__41549\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__8943\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41539\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__41539\,
            I => \N__41536\
        );

    \I__8941\ : Span4Mux_h
    port map (
            O => \N__41536\,
            I => \N__41533\
        );

    \I__8940\ : Odrv4
    port map (
            O => \N__41533\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_18\
        );

    \I__8939\ : InMux
    port map (
            O => \N__41530\,
            I => \N__41527\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__41527\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIOTCPZ0Z_18\
        );

    \I__8937\ : CascadeMux
    port map (
            O => \N__41524\,
            I => \N__41520\
        );

    \I__8936\ : InMux
    port map (
            O => \N__41523\,
            I => \N__41516\
        );

    \I__8935\ : InMux
    port map (
            O => \N__41520\,
            I => \N__41509\
        );

    \I__8934\ : InMux
    port map (
            O => \N__41519\,
            I => \N__41509\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__41516\,
            I => \N__41506\
        );

    \I__8932\ : InMux
    port map (
            O => \N__41515\,
            I => \N__41501\
        );

    \I__8931\ : InMux
    port map (
            O => \N__41514\,
            I => \N__41501\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__41509\,
            I => \N__41498\
        );

    \I__8929\ : Span4Mux_v
    port map (
            O => \N__41506\,
            I => \N__41495\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__41501\,
            I => \N__41492\
        );

    \I__8927\ : Span4Mux_h
    port map (
            O => \N__41498\,
            I => \N__41489\
        );

    \I__8926\ : Odrv4
    port map (
            O => \N__41495\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__8925\ : Odrv4
    port map (
            O => \N__41492\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__8924\ : Odrv4
    port map (
            O => \N__41489\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__8923\ : CascadeMux
    port map (
            O => \N__41482\,
            I => \N__41479\
        );

    \I__8922\ : InMux
    port map (
            O => \N__41479\,
            I => \N__41476\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__41476\,
            I => \current_shift_inst.PI_CTRL.integrator_i_14\
        );

    \I__8920\ : CascadeMux
    port map (
            O => \N__41473\,
            I => \N__41470\
        );

    \I__8919\ : InMux
    port map (
            O => \N__41470\,
            I => \N__41467\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__41467\,
            I => \current_shift_inst.PI_CTRL.integrator_i_8\
        );

    \I__8917\ : InMux
    port map (
            O => \N__41464\,
            I => \N__41461\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__41461\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__8915\ : InMux
    port map (
            O => \N__41458\,
            I => \N__41455\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__41455\,
            I => \N__41450\
        );

    \I__8913\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41447\
        );

    \I__8912\ : CascadeMux
    port map (
            O => \N__41453\,
            I => \N__41443\
        );

    \I__8911\ : Span4Mux_v
    port map (
            O => \N__41450\,
            I => \N__41438\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__41447\,
            I => \N__41438\
        );

    \I__8909\ : InMux
    port map (
            O => \N__41446\,
            I => \N__41435\
        );

    \I__8908\ : InMux
    port map (
            O => \N__41443\,
            I => \N__41432\
        );

    \I__8907\ : Span4Mux_h
    port map (
            O => \N__41438\,
            I => \N__41429\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__41435\,
            I => \N__41425\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__41432\,
            I => \N__41420\
        );

    \I__8904\ : Span4Mux_h
    port map (
            O => \N__41429\,
            I => \N__41420\
        );

    \I__8903\ : InMux
    port map (
            O => \N__41428\,
            I => \N__41417\
        );

    \I__8902\ : Odrv12
    port map (
            O => \N__41425\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__8901\ : Odrv4
    port map (
            O => \N__41420\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__41417\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__8899\ : InMux
    port map (
            O => \N__41410\,
            I => \N__41407\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__41407\,
            I => \N__41404\
        );

    \I__8897\ : Span4Mux_v
    port map (
            O => \N__41404\,
            I => \N__41401\
        );

    \I__8896\ : Odrv4
    port map (
            O => \N__41401\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_25\
        );

    \I__8895\ : InMux
    port map (
            O => \N__41398\,
            I => \N__41395\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__41395\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIGNFQZ0Z_25\
        );

    \I__8893\ : InMux
    port map (
            O => \N__41392\,
            I => \N__41387\
        );

    \I__8892\ : InMux
    port map (
            O => \N__41391\,
            I => \N__41382\
        );

    \I__8891\ : InMux
    port map (
            O => \N__41390\,
            I => \N__41382\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__41387\,
            I => \N__41379\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__41382\,
            I => \N__41376\
        );

    \I__8888\ : Span4Mux_h
    port map (
            O => \N__41379\,
            I => \N__41373\
        );

    \I__8887\ : Span4Mux_h
    port map (
            O => \N__41376\,
            I => \N__41370\
        );

    \I__8886\ : Odrv4
    port map (
            O => \N__41373\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__8885\ : Odrv4
    port map (
            O => \N__41370\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__8884\ : InMux
    port map (
            O => \N__41365\,
            I => \N__41362\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__41362\,
            I => \N__41359\
        );

    \I__8882\ : Span4Mux_h
    port map (
            O => \N__41359\,
            I => \N__41356\
        );

    \I__8881\ : Odrv4
    port map (
            O => \N__41356\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__8880\ : InMux
    port map (
            O => \N__41353\,
            I => \N__41350\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__41350\,
            I => \N__41347\
        );

    \I__8878\ : Odrv4
    port map (
            O => \N__41347\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__8877\ : InMux
    port map (
            O => \N__41344\,
            I => \N__41341\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__41341\,
            I => \N__41335\
        );

    \I__8875\ : InMux
    port map (
            O => \N__41340\,
            I => \N__41332\
        );

    \I__8874\ : InMux
    port map (
            O => \N__41339\,
            I => \N__41329\
        );

    \I__8873\ : InMux
    port map (
            O => \N__41338\,
            I => \N__41326\
        );

    \I__8872\ : Span4Mux_v
    port map (
            O => \N__41335\,
            I => \N__41323\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__41332\,
            I => \N__41320\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__41329\,
            I => \N__41316\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__41326\,
            I => \N__41313\
        );

    \I__8868\ : Span4Mux_h
    port map (
            O => \N__41323\,
            I => \N__41308\
        );

    \I__8867\ : Span4Mux_v
    port map (
            O => \N__41320\,
            I => \N__41308\
        );

    \I__8866\ : InMux
    port map (
            O => \N__41319\,
            I => \N__41305\
        );

    \I__8865\ : Span4Mux_v
    port map (
            O => \N__41316\,
            I => \N__41302\
        );

    \I__8864\ : Span4Mux_v
    port map (
            O => \N__41313\,
            I => \N__41299\
        );

    \I__8863\ : Span4Mux_h
    port map (
            O => \N__41308\,
            I => \N__41294\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__41305\,
            I => \N__41294\
        );

    \I__8861\ : Span4Mux_h
    port map (
            O => \N__41302\,
            I => \N__41291\
        );

    \I__8860\ : Odrv4
    port map (
            O => \N__41299\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__41294\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__8858\ : Odrv4
    port map (
            O => \N__41291\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__8857\ : InMux
    port map (
            O => \N__41284\,
            I => \N__41281\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__41281\,
            I => \N__41278\
        );

    \I__8855\ : Odrv4
    port map (
            O => \N__41278\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__8854\ : InMux
    port map (
            O => \N__41275\,
            I => \N__41272\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__41272\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__8852\ : InMux
    port map (
            O => \N__41269\,
            I => \N__41266\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__41266\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__8850\ : InMux
    port map (
            O => \N__41263\,
            I => \N__41260\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__41260\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\
        );

    \I__8848\ : InMux
    port map (
            O => \N__41257\,
            I => \N__41253\
        );

    \I__8847\ : InMux
    port map (
            O => \N__41256\,
            I => \N__41250\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__41253\,
            I => measured_delay_hc_29
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__41250\,
            I => measured_delay_hc_29
        );

    \I__8844\ : InMux
    port map (
            O => \N__41245\,
            I => \N__41241\
        );

    \I__8843\ : InMux
    port map (
            O => \N__41244\,
            I => \N__41238\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__41241\,
            I => measured_delay_hc_30
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__41238\,
            I => measured_delay_hc_30
        );

    \I__8840\ : InMux
    port map (
            O => \N__41233\,
            I => \N__41229\
        );

    \I__8839\ : InMux
    port map (
            O => \N__41232\,
            I => \N__41226\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__41229\,
            I => measured_delay_hc_27
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__41226\,
            I => measured_delay_hc_27
        );

    \I__8836\ : CascadeMux
    port map (
            O => \N__41221\,
            I => \N__41216\
        );

    \I__8835\ : CascadeMux
    port map (
            O => \N__41220\,
            I => \N__41204\
        );

    \I__8834\ : CascadeMux
    port map (
            O => \N__41219\,
            I => \N__41200\
        );

    \I__8833\ : InMux
    port map (
            O => \N__41216\,
            I => \N__41188\
        );

    \I__8832\ : InMux
    port map (
            O => \N__41215\,
            I => \N__41188\
        );

    \I__8831\ : InMux
    port map (
            O => \N__41214\,
            I => \N__41188\
        );

    \I__8830\ : InMux
    port map (
            O => \N__41213\,
            I => \N__41180\
        );

    \I__8829\ : InMux
    port map (
            O => \N__41212\,
            I => \N__41177\
        );

    \I__8828\ : CascadeMux
    port map (
            O => \N__41211\,
            I => \N__41174\
        );

    \I__8827\ : CascadeMux
    port map (
            O => \N__41210\,
            I => \N__41171\
        );

    \I__8826\ : CascadeMux
    port map (
            O => \N__41209\,
            I => \N__41166\
        );

    \I__8825\ : CascadeMux
    port map (
            O => \N__41208\,
            I => \N__41163\
        );

    \I__8824\ : CascadeMux
    port map (
            O => \N__41207\,
            I => \N__41160\
        );

    \I__8823\ : InMux
    port map (
            O => \N__41204\,
            I => \N__41150\
        );

    \I__8822\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41143\
        );

    \I__8821\ : InMux
    port map (
            O => \N__41200\,
            I => \N__41143\
        );

    \I__8820\ : InMux
    port map (
            O => \N__41199\,
            I => \N__41143\
        );

    \I__8819\ : InMux
    port map (
            O => \N__41198\,
            I => \N__41134\
        );

    \I__8818\ : InMux
    port map (
            O => \N__41197\,
            I => \N__41134\
        );

    \I__8817\ : InMux
    port map (
            O => \N__41196\,
            I => \N__41134\
        );

    \I__8816\ : InMux
    port map (
            O => \N__41195\,
            I => \N__41134\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__41188\,
            I => \N__41131\
        );

    \I__8814\ : InMux
    port map (
            O => \N__41187\,
            I => \N__41128\
        );

    \I__8813\ : InMux
    port map (
            O => \N__41186\,
            I => \N__41119\
        );

    \I__8812\ : InMux
    port map (
            O => \N__41185\,
            I => \N__41119\
        );

    \I__8811\ : InMux
    port map (
            O => \N__41184\,
            I => \N__41119\
        );

    \I__8810\ : InMux
    port map (
            O => \N__41183\,
            I => \N__41119\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__41180\,
            I => \N__41114\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__41177\,
            I => \N__41114\
        );

    \I__8807\ : InMux
    port map (
            O => \N__41174\,
            I => \N__41105\
        );

    \I__8806\ : InMux
    port map (
            O => \N__41171\,
            I => \N__41105\
        );

    \I__8805\ : InMux
    port map (
            O => \N__41170\,
            I => \N__41105\
        );

    \I__8804\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41105\
        );

    \I__8803\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41094\
        );

    \I__8802\ : InMux
    port map (
            O => \N__41163\,
            I => \N__41094\
        );

    \I__8801\ : InMux
    port map (
            O => \N__41160\,
            I => \N__41094\
        );

    \I__8800\ : InMux
    port map (
            O => \N__41159\,
            I => \N__41094\
        );

    \I__8799\ : InMux
    port map (
            O => \N__41158\,
            I => \N__41094\
        );

    \I__8798\ : InMux
    port map (
            O => \N__41157\,
            I => \N__41083\
        );

    \I__8797\ : InMux
    port map (
            O => \N__41156\,
            I => \N__41083\
        );

    \I__8796\ : InMux
    port map (
            O => \N__41155\,
            I => \N__41083\
        );

    \I__8795\ : InMux
    port map (
            O => \N__41154\,
            I => \N__41083\
        );

    \I__8794\ : InMux
    port map (
            O => \N__41153\,
            I => \N__41083\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__41150\,
            I => \N__41074\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__41143\,
            I => \N__41074\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__41134\,
            I => \N__41074\
        );

    \I__8790\ : Span4Mux_h
    port map (
            O => \N__41131\,
            I => \N__41074\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__41128\,
            I => \N__41071\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__41119\,
            I => \N__41068\
        );

    \I__8787\ : Span4Mux_h
    port map (
            O => \N__41114\,
            I => \N__41065\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__41105\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__41094\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__41083\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8783\ : Odrv4
    port map (
            O => \N__41074\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8782\ : Odrv12
    port map (
            O => \N__41071\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8781\ : Odrv12
    port map (
            O => \N__41068\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8780\ : Odrv4
    port map (
            O => \N__41065\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8779\ : InMux
    port map (
            O => \N__41050\,
            I => \N__41043\
        );

    \I__8778\ : InMux
    port map (
            O => \N__41049\,
            I => \N__41025\
        );

    \I__8777\ : InMux
    port map (
            O => \N__41048\,
            I => \N__41025\
        );

    \I__8776\ : InMux
    port map (
            O => \N__41047\,
            I => \N__41025\
        );

    \I__8775\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41022\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__41043\,
            I => \N__41009\
        );

    \I__8773\ : InMux
    port map (
            O => \N__41042\,
            I => \N__41002\
        );

    \I__8772\ : InMux
    port map (
            O => \N__41041\,
            I => \N__41002\
        );

    \I__8771\ : InMux
    port map (
            O => \N__41040\,
            I => \N__41002\
        );

    \I__8770\ : InMux
    port map (
            O => \N__41039\,
            I => \N__40993\
        );

    \I__8769\ : InMux
    port map (
            O => \N__41038\,
            I => \N__40993\
        );

    \I__8768\ : InMux
    port map (
            O => \N__41037\,
            I => \N__40993\
        );

    \I__8767\ : InMux
    port map (
            O => \N__41036\,
            I => \N__40993\
        );

    \I__8766\ : InMux
    port map (
            O => \N__41035\,
            I => \N__40984\
        );

    \I__8765\ : InMux
    port map (
            O => \N__41034\,
            I => \N__40984\
        );

    \I__8764\ : InMux
    port map (
            O => \N__41033\,
            I => \N__40984\
        );

    \I__8763\ : InMux
    port map (
            O => \N__41032\,
            I => \N__40984\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__41025\,
            I => \N__40975\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__41022\,
            I => \N__40972\
        );

    \I__8760\ : InMux
    port map (
            O => \N__41021\,
            I => \N__40959\
        );

    \I__8759\ : InMux
    port map (
            O => \N__41020\,
            I => \N__40959\
        );

    \I__8758\ : InMux
    port map (
            O => \N__41019\,
            I => \N__40959\
        );

    \I__8757\ : InMux
    port map (
            O => \N__41018\,
            I => \N__40959\
        );

    \I__8756\ : InMux
    port map (
            O => \N__41017\,
            I => \N__40959\
        );

    \I__8755\ : InMux
    port map (
            O => \N__41016\,
            I => \N__40959\
        );

    \I__8754\ : InMux
    port map (
            O => \N__41015\,
            I => \N__40950\
        );

    \I__8753\ : InMux
    port map (
            O => \N__41014\,
            I => \N__40950\
        );

    \I__8752\ : InMux
    port map (
            O => \N__41013\,
            I => \N__40950\
        );

    \I__8751\ : InMux
    port map (
            O => \N__41012\,
            I => \N__40950\
        );

    \I__8750\ : Span4Mux_h
    port map (
            O => \N__41009\,
            I => \N__40947\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__41002\,
            I => \N__40944\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__40993\,
            I => \N__40939\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__40984\,
            I => \N__40939\
        );

    \I__8746\ : InMux
    port map (
            O => \N__40983\,
            I => \N__40936\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40925\
        );

    \I__8744\ : InMux
    port map (
            O => \N__40981\,
            I => \N__40925\
        );

    \I__8743\ : InMux
    port map (
            O => \N__40980\,
            I => \N__40925\
        );

    \I__8742\ : InMux
    port map (
            O => \N__40979\,
            I => \N__40925\
        );

    \I__8741\ : InMux
    port map (
            O => \N__40978\,
            I => \N__40925\
        );

    \I__8740\ : Span4Mux_h
    port map (
            O => \N__40975\,
            I => \N__40916\
        );

    \I__8739\ : Span4Mux_h
    port map (
            O => \N__40972\,
            I => \N__40916\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__40959\,
            I => \N__40916\
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__40950\,
            I => \N__40916\
        );

    \I__8736\ : Odrv4
    port map (
            O => \N__40947\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8735\ : Odrv12
    port map (
            O => \N__40944\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8734\ : Odrv12
    port map (
            O => \N__40939\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__40936\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__40925\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8731\ : Odrv4
    port map (
            O => \N__40916\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8730\ : InMux
    port map (
            O => \N__40903\,
            I => \N__40899\
        );

    \I__8729\ : InMux
    port map (
            O => \N__40902\,
            I => \N__40896\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__40899\,
            I => measured_delay_hc_28
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__40896\,
            I => measured_delay_hc_28
        );

    \I__8726\ : InMux
    port map (
            O => \N__40891\,
            I => \N__40888\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__40888\,
            I => \N__40885\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__40885\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__8723\ : InMux
    port map (
            O => \N__40882\,
            I => \N__40878\
        );

    \I__8722\ : CascadeMux
    port map (
            O => \N__40881\,
            I => \N__40874\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__40878\,
            I => \N__40870\
        );

    \I__8720\ : InMux
    port map (
            O => \N__40877\,
            I => \N__40867\
        );

    \I__8719\ : InMux
    port map (
            O => \N__40874\,
            I => \N__40864\
        );

    \I__8718\ : InMux
    port map (
            O => \N__40873\,
            I => \N__40861\
        );

    \I__8717\ : Span4Mux_v
    port map (
            O => \N__40870\,
            I => \N__40858\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__40867\,
            I => \N__40855\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__40864\,
            I => \N__40851\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__40861\,
            I => \N__40844\
        );

    \I__8713\ : Span4Mux_h
    port map (
            O => \N__40858\,
            I => \N__40844\
        );

    \I__8712\ : Span4Mux_v
    port map (
            O => \N__40855\,
            I => \N__40844\
        );

    \I__8711\ : InMux
    port map (
            O => \N__40854\,
            I => \N__40841\
        );

    \I__8710\ : Span12Mux_v
    port map (
            O => \N__40851\,
            I => \N__40838\
        );

    \I__8709\ : Span4Mux_h
    port map (
            O => \N__40844\,
            I => \N__40833\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__40841\,
            I => \N__40833\
        );

    \I__8707\ : Odrv12
    port map (
            O => \N__40838\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__8706\ : Odrv4
    port map (
            O => \N__40833\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__8705\ : CascadeMux
    port map (
            O => \N__40828\,
            I => \N__40825\
        );

    \I__8704\ : InMux
    port map (
            O => \N__40825\,
            I => \N__40822\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__40822\,
            I => \N__40819\
        );

    \I__8702\ : Span4Mux_v
    port map (
            O => \N__40819\,
            I => \N__40816\
        );

    \I__8701\ : Odrv4
    port map (
            O => \N__40816\,
            I => \current_shift_inst.PI_CTRL.integrator_i_25\
        );

    \I__8700\ : InMux
    port map (
            O => \N__40813\,
            I => \N__40810\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__40810\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\
        );

    \I__8698\ : InMux
    port map (
            O => \N__40807\,
            I => \N__40804\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__40804\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__8696\ : InMux
    port map (
            O => \N__40801\,
            I => \N__40798\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__40798\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__8694\ : InMux
    port map (
            O => \N__40795\,
            I => \N__40792\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__40792\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__8692\ : InMux
    port map (
            O => \N__40789\,
            I => \N__40786\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__40786\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__8690\ : InMux
    port map (
            O => \N__40783\,
            I => \N__40780\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__40780\,
            I => \N__40777\
        );

    \I__8688\ : Span4Mux_h
    port map (
            O => \N__40777\,
            I => \N__40773\
        );

    \I__8687\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40770\
        );

    \I__8686\ : Odrv4
    port map (
            O => \N__40773\,
            I => \current_shift_inst.un4_control_input_0_31\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__40770\,
            I => \current_shift_inst.un4_control_input_0_31\
        );

    \I__8684\ : InMux
    port map (
            O => \N__40765\,
            I => \N__40762\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__40762\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__8682\ : InMux
    port map (
            O => \N__40759\,
            I => \N__40756\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__40756\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__8680\ : InMux
    port map (
            O => \N__40753\,
            I => \N__40750\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__40750\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\
        );

    \I__8678\ : CascadeMux
    port map (
            O => \N__40747\,
            I => \N__40744\
        );

    \I__8677\ : InMux
    port map (
            O => \N__40744\,
            I => \N__40741\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__40741\,
            I => \N__40738\
        );

    \I__8675\ : Odrv4
    port map (
            O => \N__40738\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__8674\ : InMux
    port map (
            O => \N__40735\,
            I => \N__40732\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__40732\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\
        );

    \I__8672\ : InMux
    port map (
            O => \N__40729\,
            I => \N__40726\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__40726\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__8670\ : InMux
    port map (
            O => \N__40723\,
            I => \N__40720\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__40720\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\
        );

    \I__8668\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40714\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__40714\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__8666\ : CascadeMux
    port map (
            O => \N__40711\,
            I => \N__40708\
        );

    \I__8665\ : InMux
    port map (
            O => \N__40708\,
            I => \N__40705\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__40705\,
            I => \N__40702\
        );

    \I__8663\ : Odrv12
    port map (
            O => \N__40702\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__8662\ : InMux
    port map (
            O => \N__40699\,
            I => \N__40696\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__40696\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\
        );

    \I__8660\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40690\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__40690\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\
        );

    \I__8658\ : InMux
    port map (
            O => \N__40687\,
            I => \N__40684\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__40684\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\
        );

    \I__8656\ : CascadeMux
    port map (
            O => \N__40681\,
            I => \N__40678\
        );

    \I__8655\ : InMux
    port map (
            O => \N__40678\,
            I => \N__40675\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__40675\,
            I => \N__40672\
        );

    \I__8653\ : Span4Mux_h
    port map (
            O => \N__40672\,
            I => \N__40669\
        );

    \I__8652\ : Odrv4
    port map (
            O => \N__40669\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__8651\ : InMux
    port map (
            O => \N__40666\,
            I => \N__40663\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__40663\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__8649\ : InMux
    port map (
            O => \N__40660\,
            I => \N__40657\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__40657\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__8647\ : InMux
    port map (
            O => \N__40654\,
            I => \N__40651\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__40651\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__8645\ : CascadeMux
    port map (
            O => \N__40648\,
            I => \N__40645\
        );

    \I__8644\ : InMux
    port map (
            O => \N__40645\,
            I => \N__40642\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__40642\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__8642\ : InMux
    port map (
            O => \N__40639\,
            I => \N__40636\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__40636\,
            I => \N__40633\
        );

    \I__8640\ : Span4Mux_v
    port map (
            O => \N__40633\,
            I => \N__40630\
        );

    \I__8639\ : Odrv4
    port map (
            O => \N__40630\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__8638\ : InMux
    port map (
            O => \N__40627\,
            I => \N__40624\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__40624\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\
        );

    \I__8636\ : InMux
    port map (
            O => \N__40621\,
            I => \N__40618\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__40618\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\
        );

    \I__8634\ : InMux
    port map (
            O => \N__40615\,
            I => \N__40612\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__40612\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__8632\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40606\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__40606\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__8630\ : InMux
    port map (
            O => \N__40603\,
            I => \N__40600\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__40600\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__8628\ : InMux
    port map (
            O => \N__40597\,
            I => \N__40594\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__40594\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__8626\ : InMux
    port map (
            O => \N__40591\,
            I => \N__40588\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__40588\,
            I => \N__40585\
        );

    \I__8624\ : Span4Mux_h
    port map (
            O => \N__40585\,
            I => \N__40582\
        );

    \I__8623\ : Odrv4
    port map (
            O => \N__40582\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\
        );

    \I__8622\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40576\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__40576\,
            I => \N__40573\
        );

    \I__8620\ : Span4Mux_v
    port map (
            O => \N__40573\,
            I => \N__40570\
        );

    \I__8619\ : Odrv4
    port map (
            O => \N__40570\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\
        );

    \I__8618\ : InMux
    port map (
            O => \N__40567\,
            I => \N__40564\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__40564\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__8616\ : InMux
    port map (
            O => \N__40561\,
            I => \N__40558\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__40558\,
            I => \N__40555\
        );

    \I__8614\ : Odrv4
    port map (
            O => \N__40555\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\
        );

    \I__8613\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40549\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__40549\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__8611\ : InMux
    port map (
            O => \N__40546\,
            I => \N__40543\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__40543\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__8609\ : InMux
    port map (
            O => \N__40540\,
            I => \N__40537\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__40537\,
            I => \N__40534\
        );

    \I__8607\ : Odrv4
    port map (
            O => \N__40534\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__8606\ : InMux
    port map (
            O => \N__40531\,
            I => \N__40528\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__40528\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__8604\ : InMux
    port map (
            O => \N__40525\,
            I => \N__40522\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__40522\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__8602\ : InMux
    port map (
            O => \N__40519\,
            I => \N__40516\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__40516\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__8600\ : InMux
    port map (
            O => \N__40513\,
            I => \N__40510\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__40510\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__8598\ : InMux
    port map (
            O => \N__40507\,
            I => \N__40504\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__40504\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__8596\ : InMux
    port map (
            O => \N__40501\,
            I => \N__40498\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__40498\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__8594\ : InMux
    port map (
            O => \N__40495\,
            I => \N__40492\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__40492\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__8592\ : InMux
    port map (
            O => \N__40489\,
            I => \N__40486\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__40486\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__8590\ : InMux
    port map (
            O => \N__40483\,
            I => \N__40480\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__40480\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__8588\ : InMux
    port map (
            O => \N__40477\,
            I => \N__40474\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__40474\,
            I => \N__40471\
        );

    \I__8586\ : Span4Mux_v
    port map (
            O => \N__40471\,
            I => \N__40468\
        );

    \I__8585\ : Odrv4
    port map (
            O => \N__40468\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__8584\ : InMux
    port map (
            O => \N__40465\,
            I => \N__40462\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__40462\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__8582\ : InMux
    port map (
            O => \N__40459\,
            I => \N__40456\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40456\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__8580\ : InMux
    port map (
            O => \N__40453\,
            I => \N__40450\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__40450\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__8578\ : CascadeMux
    port map (
            O => \N__40447\,
            I => \N__40444\
        );

    \I__8577\ : InMux
    port map (
            O => \N__40444\,
            I => \N__40441\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__40441\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__8575\ : InMux
    port map (
            O => \N__40438\,
            I => \N__40435\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__40435\,
            I => \N__40432\
        );

    \I__8573\ : Span4Mux_h
    port map (
            O => \N__40432\,
            I => \N__40429\
        );

    \I__8572\ : Odrv4
    port map (
            O => \N__40429\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__40426\,
            I => \N__40421\
        );

    \I__8570\ : CascadeMux
    port map (
            O => \N__40425\,
            I => \N__40418\
        );

    \I__8569\ : InMux
    port map (
            O => \N__40424\,
            I => \N__40412\
        );

    \I__8568\ : InMux
    port map (
            O => \N__40421\,
            I => \N__40412\
        );

    \I__8567\ : InMux
    port map (
            O => \N__40418\,
            I => \N__40409\
        );

    \I__8566\ : CascadeMux
    port map (
            O => \N__40417\,
            I => \N__40406\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__40412\,
            I => \N__40403\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__40409\,
            I => \N__40400\
        );

    \I__8563\ : InMux
    port map (
            O => \N__40406\,
            I => \N__40397\
        );

    \I__8562\ : Span4Mux_h
    port map (
            O => \N__40403\,
            I => \N__40392\
        );

    \I__8561\ : Span4Mux_h
    port map (
            O => \N__40400\,
            I => \N__40392\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__40397\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__8559\ : Odrv4
    port map (
            O => \N__40392\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__8558\ : InMux
    port map (
            O => \N__40387\,
            I => \N__40384\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__40384\,
            I => \N__40381\
        );

    \I__8556\ : Span4Mux_v
    port map (
            O => \N__40381\,
            I => \N__40378\
        );

    \I__8555\ : Odrv4
    port map (
            O => \N__40378\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__8554\ : InMux
    port map (
            O => \N__40375\,
            I => \N__40365\
        );

    \I__8553\ : InMux
    port map (
            O => \N__40374\,
            I => \N__40365\
        );

    \I__8552\ : InMux
    port map (
            O => \N__40373\,
            I => \N__40365\
        );

    \I__8551\ : InMux
    port map (
            O => \N__40372\,
            I => \N__40362\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__40365\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__40362\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8548\ : InMux
    port map (
            O => \N__40357\,
            I => \N__40354\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__40354\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__8546\ : CascadeMux
    port map (
            O => \N__40351\,
            I => \N__40348\
        );

    \I__8545\ : InMux
    port map (
            O => \N__40348\,
            I => \N__40345\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__40345\,
            I => \N__40342\
        );

    \I__8543\ : Odrv4
    port map (
            O => \N__40342\,
            I => \current_shift_inst.PI_CTRL.integrator_i_18\
        );

    \I__8542\ : InMux
    port map (
            O => \N__40339\,
            I => \N__40336\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__40336\,
            I => \N__40333\
        );

    \I__8540\ : Odrv12
    port map (
            O => \N__40333\,
            I => \current_shift_inst.PI_CTRL.integrator_i_19\
        );

    \I__8539\ : InMux
    port map (
            O => \N__40330\,
            I => \N__40327\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__40327\,
            I => \N__40322\
        );

    \I__8537\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40319\
        );

    \I__8536\ : InMux
    port map (
            O => \N__40325\,
            I => \N__40316\
        );

    \I__8535\ : Span4Mux_h
    port map (
            O => \N__40322\,
            I => \N__40313\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__40319\,
            I => \N__40310\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__40316\,
            I => \N__40307\
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__40313\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__8531\ : Odrv4
    port map (
            O => \N__40310\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__8530\ : Odrv4
    port map (
            O => \N__40307\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__8529\ : InMux
    port map (
            O => \N__40300\,
            I => \N__40297\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__40297\,
            I => \N__40294\
        );

    \I__8527\ : Span4Mux_v
    port map (
            O => \N__40294\,
            I => \N__40291\
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__40291\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_24\
        );

    \I__8525\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40285\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__40285\,
            I => \N__40282\
        );

    \I__8523\ : Odrv4
    port map (
            O => \N__40282\,
            I => \current_shift_inst.PI_CTRL.error_control_RNICIEQZ0Z_24\
        );

    \I__8522\ : InMux
    port map (
            O => \N__40279\,
            I => \N__40276\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__40276\,
            I => \N__40273\
        );

    \I__8520\ : Odrv4
    port map (
            O => \N__40273\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__8519\ : CascadeMux
    port map (
            O => \N__40270\,
            I => \N__40266\
        );

    \I__8518\ : InMux
    port map (
            O => \N__40269\,
            I => \N__40263\
        );

    \I__8517\ : InMux
    port map (
            O => \N__40266\,
            I => \N__40260\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__40263\,
            I => \N__40255\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__40260\,
            I => \N__40252\
        );

    \I__8514\ : InMux
    port map (
            O => \N__40259\,
            I => \N__40249\
        );

    \I__8513\ : CascadeMux
    port map (
            O => \N__40258\,
            I => \N__40246\
        );

    \I__8512\ : Span4Mux_h
    port map (
            O => \N__40255\,
            I => \N__40241\
        );

    \I__8511\ : Span4Mux_v
    port map (
            O => \N__40252\,
            I => \N__40241\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__40249\,
            I => \N__40237\
        );

    \I__8509\ : InMux
    port map (
            O => \N__40246\,
            I => \N__40234\
        );

    \I__8508\ : Span4Mux_h
    port map (
            O => \N__40241\,
            I => \N__40231\
        );

    \I__8507\ : InMux
    port map (
            O => \N__40240\,
            I => \N__40228\
        );

    \I__8506\ : Span4Mux_h
    port map (
            O => \N__40237\,
            I => \N__40225\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__40234\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__8504\ : Odrv4
    port map (
            O => \N__40231\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__40228\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__8502\ : Odrv4
    port map (
            O => \N__40225\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__8501\ : InMux
    port map (
            O => \N__40216\,
            I => \N__40213\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__40213\,
            I => \N__40210\
        );

    \I__8499\ : Odrv4
    port map (
            O => \N__40210\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__8498\ : CascadeMux
    port map (
            O => \N__40207\,
            I => \N__40202\
        );

    \I__8497\ : InMux
    port map (
            O => \N__40206\,
            I => \N__40199\
        );

    \I__8496\ : InMux
    port map (
            O => \N__40205\,
            I => \N__40196\
        );

    \I__8495\ : InMux
    port map (
            O => \N__40202\,
            I => \N__40192\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__40199\,
            I => \N__40189\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__40196\,
            I => \N__40186\
        );

    \I__8492\ : InMux
    port map (
            O => \N__40195\,
            I => \N__40183\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__40192\,
            I => \N__40179\
        );

    \I__8490\ : Span4Mux_h
    port map (
            O => \N__40189\,
            I => \N__40172\
        );

    \I__8489\ : Span4Mux_v
    port map (
            O => \N__40186\,
            I => \N__40172\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__40183\,
            I => \N__40172\
        );

    \I__8487\ : InMux
    port map (
            O => \N__40182\,
            I => \N__40169\
        );

    \I__8486\ : Span4Mux_v
    port map (
            O => \N__40179\,
            I => \N__40164\
        );

    \I__8485\ : Span4Mux_h
    port map (
            O => \N__40172\,
            I => \N__40164\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__40169\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__8483\ : Odrv4
    port map (
            O => \N__40164\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__8482\ : InMux
    port map (
            O => \N__40159\,
            I => \N__40156\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__40156\,
            I => \N__40153\
        );

    \I__8480\ : Odrv4
    port map (
            O => \N__40153\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__8479\ : CascadeMux
    port map (
            O => \N__40150\,
            I => \N__40146\
        );

    \I__8478\ : InMux
    port map (
            O => \N__40149\,
            I => \N__40143\
        );

    \I__8477\ : InMux
    port map (
            O => \N__40146\,
            I => \N__40138\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__40143\,
            I => \N__40135\
        );

    \I__8475\ : InMux
    port map (
            O => \N__40142\,
            I => \N__40132\
        );

    \I__8474\ : InMux
    port map (
            O => \N__40141\,
            I => \N__40129\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__40138\,
            I => \N__40126\
        );

    \I__8472\ : Span4Mux_v
    port map (
            O => \N__40135\,
            I => \N__40123\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__40132\,
            I => \N__40118\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__40129\,
            I => \N__40118\
        );

    \I__8469\ : Span4Mux_v
    port map (
            O => \N__40126\,
            I => \N__40114\
        );

    \I__8468\ : Span4Mux_h
    port map (
            O => \N__40123\,
            I => \N__40109\
        );

    \I__8467\ : Span4Mux_v
    port map (
            O => \N__40118\,
            I => \N__40109\
        );

    \I__8466\ : InMux
    port map (
            O => \N__40117\,
            I => \N__40106\
        );

    \I__8465\ : Odrv4
    port map (
            O => \N__40114\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__8464\ : Odrv4
    port map (
            O => \N__40109\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__40106\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__8462\ : InMux
    port map (
            O => \N__40099\,
            I => \N__40096\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__40096\,
            I => \N__40093\
        );

    \I__8460\ : Span4Mux_h
    port map (
            O => \N__40093\,
            I => \N__40090\
        );

    \I__8459\ : Odrv4
    port map (
            O => \N__40090\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__8458\ : InMux
    port map (
            O => \N__40087\,
            I => \N__40084\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__40084\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJZ0\
        );

    \I__8456\ : InMux
    port map (
            O => \N__40081\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\
        );

    \I__8455\ : InMux
    port map (
            O => \N__40078\,
            I => \N__40075\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__40075\,
            I => \N__40072\
        );

    \I__8453\ : Span4Mux_h
    port map (
            O => \N__40072\,
            I => \N__40069\
        );

    \I__8452\ : Odrv4
    port map (
            O => \N__40069\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5KZ0\
        );

    \I__8451\ : CascadeMux
    port map (
            O => \N__40066\,
            I => \N__40063\
        );

    \I__8450\ : InMux
    port map (
            O => \N__40063\,
            I => \N__40060\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__40060\,
            I => \N__40057\
        );

    \I__8448\ : Odrv4
    port map (
            O => \N__40057\,
            I => \current_shift_inst.PI_CTRL.integrator_i_27\
        );

    \I__8447\ : InMux
    port map (
            O => \N__40054\,
            I => \N__40051\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__40051\,
            I => \N__40048\
        );

    \I__8445\ : Odrv12
    port map (
            O => \N__40048\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__8444\ : InMux
    port map (
            O => \N__40045\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\
        );

    \I__8443\ : InMux
    port map (
            O => \N__40042\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\
        );

    \I__8442\ : InMux
    port map (
            O => \N__40039\,
            I => \N__40036\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__40036\,
            I => \N__40033\
        );

    \I__8440\ : Odrv12
    port map (
            O => \N__40033\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__8439\ : InMux
    port map (
            O => \N__40030\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\
        );

    \I__8438\ : CascadeMux
    port map (
            O => \N__40027\,
            I => \N__40024\
        );

    \I__8437\ : InMux
    port map (
            O => \N__40024\,
            I => \N__40021\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__40021\,
            I => \N__40018\
        );

    \I__8435\ : Span4Mux_h
    port map (
            O => \N__40018\,
            I => \N__40015\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__40015\,
            I => \current_shift_inst.PI_CTRL.integrator_i_30\
        );

    \I__8433\ : InMux
    port map (
            O => \N__40012\,
            I => \N__40009\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__40009\,
            I => \N__40006\
        );

    \I__8431\ : Odrv12
    port map (
            O => \N__40006\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__8430\ : InMux
    port map (
            O => \N__40003\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\
        );

    \I__8429\ : InMux
    port map (
            O => \N__40000\,
            I => \bfn_16_12_0_\
        );

    \I__8428\ : InMux
    port map (
            O => \N__39997\,
            I => \N__39993\
        );

    \I__8427\ : CascadeMux
    port map (
            O => \N__39996\,
            I => \N__39990\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__39993\,
            I => \N__39986\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39990\,
            I => \N__39982\
        );

    \I__8424\ : InMux
    port map (
            O => \N__39989\,
            I => \N__39979\
        );

    \I__8423\ : Span4Mux_h
    port map (
            O => \N__39986\,
            I => \N__39976\
        );

    \I__8422\ : InMux
    port map (
            O => \N__39985\,
            I => \N__39973\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__39982\,
            I => \N__39970\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__39979\,
            I => \N__39963\
        );

    \I__8419\ : Span4Mux_h
    port map (
            O => \N__39976\,
            I => \N__39963\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__39973\,
            I => \N__39963\
        );

    \I__8417\ : Odrv4
    port map (
            O => \N__39970\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__8416\ : Odrv4
    port map (
            O => \N__39963\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__8415\ : InMux
    port map (
            O => \N__39958\,
            I => \N__39955\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__39955\,
            I => \current_shift_inst.PI_CTRL.integrator_i_29\
        );

    \I__8413\ : CascadeMux
    port map (
            O => \N__39952\,
            I => \N__39949\
        );

    \I__8412\ : InMux
    port map (
            O => \N__39949\,
            I => \N__39946\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__39946\,
            I => \N__39943\
        );

    \I__8410\ : Odrv4
    port map (
            O => \N__39943\,
            I => \current_shift_inst.PI_CTRL.integrator_i_20\
        );

    \I__8409\ : CascadeMux
    port map (
            O => \N__39940\,
            I => \N__39936\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39939\,
            I => \N__39928\
        );

    \I__8407\ : InMux
    port map (
            O => \N__39936\,
            I => \N__39928\
        );

    \I__8406\ : InMux
    port map (
            O => \N__39935\,
            I => \N__39928\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__39928\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_0_26\
        );

    \I__8404\ : InMux
    port map (
            O => \N__39925\,
            I => \N__39922\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__39922\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIDGBQZ0Z_22\
        );

    \I__8402\ : InMux
    port map (
            O => \N__39919\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\
        );

    \I__8401\ : CascadeMux
    port map (
            O => \N__39916\,
            I => \N__39913\
        );

    \I__8400\ : InMux
    port map (
            O => \N__39913\,
            I => \N__39910\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__39910\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIHLCQZ0Z_23\
        );

    \I__8398\ : InMux
    port map (
            O => \N__39907\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\
        );

    \I__8397\ : InMux
    port map (
            O => \N__39904\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\
        );

    \I__8396\ : CascadeMux
    port map (
            O => \N__39901\,
            I => \N__39898\
        );

    \I__8395\ : InMux
    port map (
            O => \N__39898\,
            I => \N__39895\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__39895\,
            I => \N__39892\
        );

    \I__8393\ : Span4Mux_v
    port map (
            O => \N__39892\,
            I => \N__39889\
        );

    \I__8392\ : Odrv4
    port map (
            O => \N__39889\,
            I => \current_shift_inst.PI_CTRL.integrator_i_21\
        );

    \I__8391\ : InMux
    port map (
            O => \N__39886\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\
        );

    \I__8390\ : InMux
    port map (
            O => \N__39883\,
            I => \N__39880\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__39880\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7JZ0\
        );

    \I__8388\ : CascadeMux
    port map (
            O => \N__39877\,
            I => \N__39874\
        );

    \I__8387\ : InMux
    port map (
            O => \N__39874\,
            I => \N__39871\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__39871\,
            I => \N__39868\
        );

    \I__8385\ : Span4Mux_v
    port map (
            O => \N__39868\,
            I => \N__39865\
        );

    \I__8384\ : Odrv4
    port map (
            O => \N__39865\,
            I => \current_shift_inst.PI_CTRL.integrator_i_22\
        );

    \I__8383\ : InMux
    port map (
            O => \N__39862\,
            I => \N__39859\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__39859\,
            I => \N__39856\
        );

    \I__8381\ : Odrv12
    port map (
            O => \N__39856\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__8380\ : InMux
    port map (
            O => \N__39853\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\
        );

    \I__8379\ : InMux
    port map (
            O => \N__39850\,
            I => \N__39847\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__39847\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8JZ0\
        );

    \I__8377\ : InMux
    port map (
            O => \N__39844\,
            I => \bfn_16_11_0_\
        );

    \I__8376\ : InMux
    port map (
            O => \N__39841\,
            I => \N__39838\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__39838\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9JZ0\
        );

    \I__8374\ : InMux
    port map (
            O => \N__39835\,
            I => \N__39832\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__39832\,
            I => \N__39829\
        );

    \I__8372\ : Odrv12
    port map (
            O => \N__39829\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__8371\ : InMux
    port map (
            O => \N__39826\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\
        );

    \I__8370\ : InMux
    port map (
            O => \N__39823\,
            I => \N__39820\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__39820\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJZ0\
        );

    \I__8368\ : InMux
    port map (
            O => \N__39817\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\
        );

    \I__8367\ : InMux
    port map (
            O => \N__39814\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\
        );

    \I__8366\ : InMux
    port map (
            O => \N__39811\,
            I => \N__39808\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__39808\,
            I => \current_shift_inst.PI_CTRL.error_control_RNICE9PZ0Z_15\
        );

    \I__8364\ : CascadeMux
    port map (
            O => \N__39805\,
            I => \N__39802\
        );

    \I__8363\ : InMux
    port map (
            O => \N__39802\,
            I => \N__39799\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__39799\,
            I => \current_shift_inst.PI_CTRL.integrator_i_11\
        );

    \I__8361\ : InMux
    port map (
            O => \N__39796\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\
        );

    \I__8360\ : InMux
    port map (
            O => \N__39793\,
            I => \N__39790\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__39790\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIGJAPZ0Z_16\
        );

    \I__8358\ : InMux
    port map (
            O => \N__39787\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\
        );

    \I__8357\ : InMux
    port map (
            O => \N__39784\,
            I => \N__39781\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__39781\,
            I => \N__39778\
        );

    \I__8355\ : Span4Mux_h
    port map (
            O => \N__39778\,
            I => \N__39775\
        );

    \I__8354\ : Odrv4
    port map (
            O => \N__39775\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__8353\ : InMux
    port map (
            O => \N__39772\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\
        );

    \I__8352\ : InMux
    port map (
            O => \N__39769\,
            I => \N__39766\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__39766\,
            I => \N__39763\
        );

    \I__8350\ : Span4Mux_h
    port map (
            O => \N__39763\,
            I => \N__39760\
        );

    \I__8349\ : Odrv4
    port map (
            O => \N__39760\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__8348\ : InMux
    port map (
            O => \N__39757\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\
        );

    \I__8347\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39751\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__39751\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIS2EPZ0Z_19\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__39748\,
            I => \N__39745\
        );

    \I__8344\ : InMux
    port map (
            O => \N__39745\,
            I => \N__39742\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__39742\,
            I => \N__39739\
        );

    \I__8342\ : Odrv12
    port map (
            O => \N__39739\,
            I => \current_shift_inst.PI_CTRL.integrator_i_15\
        );

    \I__8341\ : InMux
    port map (
            O => \N__39736\,
            I => \N__39733\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__39733\,
            I => \N__39730\
        );

    \I__8339\ : Span4Mux_h
    port map (
            O => \N__39730\,
            I => \N__39727\
        );

    \I__8338\ : Odrv4
    port map (
            O => \N__39727\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__8337\ : InMux
    port map (
            O => \N__39724\,
            I => \bfn_16_10_0_\
        );

    \I__8336\ : InMux
    port map (
            O => \N__39721\,
            I => \N__39718\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__39718\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIENGPZ0Z_20\
        );

    \I__8334\ : CascadeMux
    port map (
            O => \N__39715\,
            I => \N__39712\
        );

    \I__8333\ : InMux
    port map (
            O => \N__39712\,
            I => \N__39709\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__39709\,
            I => \current_shift_inst.PI_CTRL.integrator_i_16\
        );

    \I__8331\ : InMux
    port map (
            O => \N__39706\,
            I => \N__39703\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__39703\,
            I => \N__39700\
        );

    \I__8329\ : Span4Mux_h
    port map (
            O => \N__39700\,
            I => \N__39697\
        );

    \I__8328\ : Odrv4
    port map (
            O => \N__39697\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__8327\ : InMux
    port map (
            O => \N__39694\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\
        );

    \I__8326\ : CascadeMux
    port map (
            O => \N__39691\,
            I => \N__39688\
        );

    \I__8325\ : InMux
    port map (
            O => \N__39688\,
            I => \N__39685\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__39685\,
            I => \N__39682\
        );

    \I__8323\ : Span4Mux_v
    port map (
            O => \N__39682\,
            I => \N__39679\
        );

    \I__8322\ : Odrv4
    port map (
            O => \N__39679\,
            I => \current_shift_inst.PI_CTRL.integrator_i_17\
        );

    \I__8321\ : InMux
    port map (
            O => \N__39676\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\
        );

    \I__8320\ : InMux
    port map (
            O => \N__39673\,
            I => \N__39670\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__39670\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIC46UZ0Z_6\
        );

    \I__8318\ : CascadeMux
    port map (
            O => \N__39667\,
            I => \N__39664\
        );

    \I__8317\ : InMux
    port map (
            O => \N__39664\,
            I => \N__39661\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__39661\,
            I => \current_shift_inst.PI_CTRL.integrator_i_2\
        );

    \I__8315\ : InMux
    port map (
            O => \N__39658\,
            I => \N__39655\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__39655\,
            I => \N__39652\
        );

    \I__8313\ : Odrv4
    port map (
            O => \N__39652\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__8312\ : InMux
    port map (
            O => \N__39649\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\
        );

    \I__8311\ : InMux
    port map (
            O => \N__39646\,
            I => \N__39643\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__39643\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIG97UZ0Z_7\
        );

    \I__8309\ : CascadeMux
    port map (
            O => \N__39640\,
            I => \N__39637\
        );

    \I__8308\ : InMux
    port map (
            O => \N__39637\,
            I => \N__39634\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__39634\,
            I => \current_shift_inst.PI_CTRL.integrator_i_3\
        );

    \I__8306\ : InMux
    port map (
            O => \N__39631\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\
        );

    \I__8305\ : InMux
    port map (
            O => \N__39628\,
            I => \N__39625\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__39625\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIKE8UZ0Z_8\
        );

    \I__8303\ : CascadeMux
    port map (
            O => \N__39622\,
            I => \N__39619\
        );

    \I__8302\ : InMux
    port map (
            O => \N__39619\,
            I => \N__39616\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__39616\,
            I => \current_shift_inst.PI_CTRL.integrator_i_4\
        );

    \I__8300\ : InMux
    port map (
            O => \N__39613\,
            I => \N__39610\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__39610\,
            I => \N__39607\
        );

    \I__8298\ : Odrv4
    port map (
            O => \N__39607\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__8297\ : InMux
    port map (
            O => \N__39604\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\
        );

    \I__8296\ : InMux
    port map (
            O => \N__39601\,
            I => \N__39598\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__39598\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIOJ9UZ0Z_9\
        );

    \I__8294\ : CascadeMux
    port map (
            O => \N__39595\,
            I => \N__39592\
        );

    \I__8293\ : InMux
    port map (
            O => \N__39592\,
            I => \N__39589\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__39589\,
            I => \N__39586\
        );

    \I__8291\ : Span4Mux_h
    port map (
            O => \N__39586\,
            I => \N__39583\
        );

    \I__8290\ : Odrv4
    port map (
            O => \N__39583\,
            I => \current_shift_inst.PI_CTRL.integrator_i_5\
        );

    \I__8289\ : InMux
    port map (
            O => \N__39580\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\
        );

    \I__8288\ : InMux
    port map (
            O => \N__39577\,
            I => \N__39574\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__39574\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIA1B41Z0Z_10\
        );

    \I__8286\ : CascadeMux
    port map (
            O => \N__39571\,
            I => \N__39568\
        );

    \I__8285\ : InMux
    port map (
            O => \N__39568\,
            I => \N__39565\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__39565\,
            I => \current_shift_inst.PI_CTRL.integrator_i_6\
        );

    \I__8283\ : InMux
    port map (
            O => \N__39562\,
            I => \N__39559\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__39559\,
            I => \N__39556\
        );

    \I__8281\ : Odrv12
    port map (
            O => \N__39556\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__8280\ : InMux
    port map (
            O => \N__39553\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\
        );

    \I__8279\ : InMux
    port map (
            O => \N__39550\,
            I => \N__39547\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__39547\,
            I => \N__39544\
        );

    \I__8277\ : Odrv4
    port map (
            O => \N__39544\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIL0S01Z0Z_11\
        );

    \I__8276\ : InMux
    port map (
            O => \N__39541\,
            I => \bfn_16_9_0_\
        );

    \I__8275\ : InMux
    port map (
            O => \N__39538\,
            I => \N__39535\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__39535\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIP5T01Z0Z_12\
        );

    \I__8273\ : InMux
    port map (
            O => \N__39532\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\
        );

    \I__8272\ : InMux
    port map (
            O => \N__39529\,
            I => \N__39526\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__39526\,
            I => \N__39523\
        );

    \I__8270\ : Span4Mux_v
    port map (
            O => \N__39523\,
            I => \N__39520\
        );

    \I__8269\ : Odrv4
    port map (
            O => \N__39520\,
            I => \current_shift_inst.PI_CTRL.error_control_RNITAU01Z0Z_13\
        );

    \I__8268\ : CascadeMux
    port map (
            O => \N__39517\,
            I => \N__39514\
        );

    \I__8267\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39511\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__39511\,
            I => \N__39508\
        );

    \I__8265\ : Odrv4
    port map (
            O => \N__39508\,
            I => \current_shift_inst.PI_CTRL.integrator_i_9\
        );

    \I__8264\ : InMux
    port map (
            O => \N__39505\,
            I => \N__39502\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__39502\,
            I => \N__39499\
        );

    \I__8262\ : Odrv4
    port map (
            O => \N__39499\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__8261\ : InMux
    port map (
            O => \N__39496\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\
        );

    \I__8260\ : CascadeMux
    port map (
            O => \N__39493\,
            I => \N__39488\
        );

    \I__8259\ : CascadeMux
    port map (
            O => \N__39492\,
            I => \N__39485\
        );

    \I__8258\ : InMux
    port map (
            O => \N__39491\,
            I => \N__39482\
        );

    \I__8257\ : InMux
    port map (
            O => \N__39488\,
            I => \N__39479\
        );

    \I__8256\ : InMux
    port map (
            O => \N__39485\,
            I => \N__39475\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__39482\,
            I => \N__39472\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__39479\,
            I => \N__39469\
        );

    \I__8253\ : InMux
    port map (
            O => \N__39478\,
            I => \N__39466\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__39475\,
            I => \N__39462\
        );

    \I__8251\ : Span4Mux_h
    port map (
            O => \N__39472\,
            I => \N__39455\
        );

    \I__8250\ : Span4Mux_v
    port map (
            O => \N__39469\,
            I => \N__39455\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__39466\,
            I => \N__39455\
        );

    \I__8248\ : InMux
    port map (
            O => \N__39465\,
            I => \N__39452\
        );

    \I__8247\ : Span4Mux_v
    port map (
            O => \N__39462\,
            I => \N__39449\
        );

    \I__8246\ : Span4Mux_v
    port map (
            O => \N__39455\,
            I => \N__39446\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__39452\,
            I => \N__39443\
        );

    \I__8244\ : Odrv4
    port map (
            O => \N__39449\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__8243\ : Odrv4
    port map (
            O => \N__39446\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__8242\ : Odrv4
    port map (
            O => \N__39443\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__8241\ : InMux
    port map (
            O => \N__39436\,
            I => \N__39433\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__39433\,
            I => \N__39429\
        );

    \I__8239\ : InMux
    port map (
            O => \N__39432\,
            I => \N__39426\
        );

    \I__8238\ : Span4Mux_v
    port map (
            O => \N__39429\,
            I => \N__39422\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__39426\,
            I => \N__39419\
        );

    \I__8236\ : InMux
    port map (
            O => \N__39425\,
            I => \N__39416\
        );

    \I__8235\ : Span4Mux_h
    port map (
            O => \N__39422\,
            I => \N__39413\
        );

    \I__8234\ : Span4Mux_h
    port map (
            O => \N__39419\,
            I => \N__39408\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__39416\,
            I => \N__39408\
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__39413\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__8231\ : Odrv4
    port map (
            O => \N__39408\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__8230\ : CascadeMux
    port map (
            O => \N__39403\,
            I => \N__39399\
        );

    \I__8229\ : InMux
    port map (
            O => \N__39402\,
            I => \N__39396\
        );

    \I__8228\ : InMux
    port map (
            O => \N__39399\,
            I => \N__39393\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__39396\,
            I => \N__39389\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__39393\,
            I => \N__39386\
        );

    \I__8225\ : CascadeMux
    port map (
            O => \N__39392\,
            I => \N__39383\
        );

    \I__8224\ : Span4Mux_v
    port map (
            O => \N__39389\,
            I => \N__39378\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__39386\,
            I => \N__39378\
        );

    \I__8222\ : InMux
    port map (
            O => \N__39383\,
            I => \N__39374\
        );

    \I__8221\ : Span4Mux_h
    port map (
            O => \N__39378\,
            I => \N__39371\
        );

    \I__8220\ : InMux
    port map (
            O => \N__39377\,
            I => \N__39368\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__39374\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__8218\ : Odrv4
    port map (
            O => \N__39371\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__39368\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__8216\ : CascadeMux
    port map (
            O => \N__39361\,
            I => \N__39357\
        );

    \I__8215\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39354\
        );

    \I__8214\ : InMux
    port map (
            O => \N__39357\,
            I => \N__39350\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__39354\,
            I => \N__39347\
        );

    \I__8212\ : InMux
    port map (
            O => \N__39353\,
            I => \N__39344\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__39350\,
            I => \N__39338\
        );

    \I__8210\ : Span4Mux_h
    port map (
            O => \N__39347\,
            I => \N__39338\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__39344\,
            I => \N__39335\
        );

    \I__8208\ : InMux
    port map (
            O => \N__39343\,
            I => \N__39332\
        );

    \I__8207\ : Span4Mux_h
    port map (
            O => \N__39338\,
            I => \N__39328\
        );

    \I__8206\ : Span4Mux_h
    port map (
            O => \N__39335\,
            I => \N__39325\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__39332\,
            I => \N__39322\
        );

    \I__8204\ : InMux
    port map (
            O => \N__39331\,
            I => \N__39319\
        );

    \I__8203\ : Odrv4
    port map (
            O => \N__39328\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__8202\ : Odrv4
    port map (
            O => \N__39325\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__8201\ : Odrv12
    port map (
            O => \N__39322\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__39319\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__8199\ : CascadeMux
    port map (
            O => \N__39310\,
            I => \N__39306\
        );

    \I__8198\ : InMux
    port map (
            O => \N__39309\,
            I => \N__39303\
        );

    \I__8197\ : InMux
    port map (
            O => \N__39306\,
            I => \N__39300\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__39303\,
            I => \N__39297\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__39300\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_26\
        );

    \I__8194\ : Odrv4
    port map (
            O => \N__39297\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_26\
        );

    \I__8193\ : InMux
    port map (
            O => \N__39292\,
            I => \N__39289\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__39289\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI4Q3UZ0Z_4\
        );

    \I__8191\ : CascadeMux
    port map (
            O => \N__39286\,
            I => \N__39282\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__39285\,
            I => \N__39279\
        );

    \I__8189\ : InMux
    port map (
            O => \N__39282\,
            I => \N__39276\
        );

    \I__8188\ : InMux
    port map (
            O => \N__39279\,
            I => \N__39273\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__39276\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__39273\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__8185\ : InMux
    port map (
            O => \N__39268\,
            I => \N__39265\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__39265\,
            I => \N__39262\
        );

    \I__8183\ : Odrv4
    port map (
            O => \N__39262\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\
        );

    \I__8182\ : InMux
    port map (
            O => \N__39259\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\
        );

    \I__8181\ : InMux
    port map (
            O => \N__39256\,
            I => \N__39253\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__39253\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI8V4UZ0Z_5\
        );

    \I__8179\ : CascadeMux
    port map (
            O => \N__39250\,
            I => \N__39247\
        );

    \I__8178\ : InMux
    port map (
            O => \N__39247\,
            I => \N__39244\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__39244\,
            I => \current_shift_inst.PI_CTRL.integrator_i_1\
        );

    \I__8176\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39238\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__39238\,
            I => \N__39235\
        );

    \I__8174\ : Span4Mux_h
    port map (
            O => \N__39235\,
            I => \N__39232\
        );

    \I__8173\ : Span4Mux_h
    port map (
            O => \N__39232\,
            I => \N__39229\
        );

    \I__8172\ : Odrv4
    port map (
            O => \N__39229\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\
        );

    \I__8171\ : InMux
    port map (
            O => \N__39226\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\
        );

    \I__8170\ : IoInMux
    port map (
            O => \N__39223\,
            I => \N__39220\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__39220\,
            I => \N__39217\
        );

    \I__8168\ : Span4Mux_s1_v
    port map (
            O => \N__39217\,
            I => \N__39214\
        );

    \I__8167\ : Span4Mux_h
    port map (
            O => \N__39214\,
            I => \N__39211\
        );

    \I__8166\ : Odrv4
    port map (
            O => \N__39211\,
            I => \delay_measurement_inst.delay_tr_timer.N_304_i\
        );

    \I__8165\ : InMux
    port map (
            O => \N__39208\,
            I => \N__39203\
        );

    \I__8164\ : InMux
    port map (
            O => \N__39207\,
            I => \N__39200\
        );

    \I__8163\ : InMux
    port map (
            O => \N__39206\,
            I => \N__39197\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__39203\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__39200\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__39197\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__8159\ : InMux
    port map (
            O => \N__39190\,
            I => \N__39182\
        );

    \I__8158\ : InMux
    port map (
            O => \N__39189\,
            I => \N__39182\
        );

    \I__8157\ : InMux
    port map (
            O => \N__39188\,
            I => \N__39179\
        );

    \I__8156\ : InMux
    port map (
            O => \N__39187\,
            I => \N__39176\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__39182\,
            I => delay_tr_d2
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__39179\,
            I => delay_tr_d2
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__39176\,
            I => delay_tr_d2
        );

    \I__8152\ : InMux
    port map (
            O => \N__39169\,
            I => \N__39164\
        );

    \I__8151\ : InMux
    port map (
            O => \N__39168\,
            I => \N__39161\
        );

    \I__8150\ : InMux
    port map (
            O => \N__39167\,
            I => \N__39158\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__39164\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__39161\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__39158\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__8146\ : InMux
    port map (
            O => \N__39151\,
            I => \N__39147\
        );

    \I__8145\ : InMux
    port map (
            O => \N__39150\,
            I => \N__39144\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__39147\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__39144\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__8142\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39135\
        );

    \I__8141\ : InMux
    port map (
            O => \N__39138\,
            I => \N__39131\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__39135\,
            I => \N__39128\
        );

    \I__8139\ : InMux
    port map (
            O => \N__39134\,
            I => \N__39125\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__39131\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__8137\ : Odrv4
    port map (
            O => \N__39128\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__39125\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__8135\ : InMux
    port map (
            O => \N__39118\,
            I => \N__39112\
        );

    \I__8134\ : InMux
    port map (
            O => \N__39117\,
            I => \N__39107\
        );

    \I__8133\ : InMux
    port map (
            O => \N__39116\,
            I => \N__39107\
        );

    \I__8132\ : InMux
    port map (
            O => \N__39115\,
            I => \N__39104\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__39112\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__39107\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__39104\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8128\ : InMux
    port map (
            O => \N__39097\,
            I => \N__39094\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__39094\,
            I => \N__39091\
        );

    \I__8126\ : Span4Mux_h
    port map (
            O => \N__39091\,
            I => \N__39088\
        );

    \I__8125\ : Odrv4
    port map (
            O => \N__39088\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__8124\ : InMux
    port map (
            O => \N__39085\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__8123\ : InMux
    port map (
            O => \N__39082\,
            I => \N__39079\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__39079\,
            I => \N__39076\
        );

    \I__8121\ : Span4Mux_v
    port map (
            O => \N__39076\,
            I => \N__39073\
        );

    \I__8120\ : Odrv4
    port map (
            O => \N__39073\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__8119\ : InMux
    port map (
            O => \N__39070\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__8118\ : InMux
    port map (
            O => \N__39067\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__8117\ : InMux
    port map (
            O => \N__39064\,
            I => \N__39061\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__39061\,
            I => \N__39058\
        );

    \I__8115\ : Span4Mux_h
    port map (
            O => \N__39058\,
            I => \N__39055\
        );

    \I__8114\ : Odrv4
    port map (
            O => \N__39055\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__8113\ : InMux
    port map (
            O => \N__39052\,
            I => \N__39049\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__39049\,
            I => \N__39044\
        );

    \I__8111\ : InMux
    port map (
            O => \N__39048\,
            I => \N__39041\
        );

    \I__8110\ : CascadeMux
    port map (
            O => \N__39047\,
            I => \N__39038\
        );

    \I__8109\ : Span4Mux_h
    port map (
            O => \N__39044\,
            I => \N__39035\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__39041\,
            I => \N__39032\
        );

    \I__8107\ : InMux
    port map (
            O => \N__39038\,
            I => \N__39029\
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__39035\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__8105\ : Odrv4
    port map (
            O => \N__39032\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__39029\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__8103\ : InMux
    port map (
            O => \N__39022\,
            I => \N__39019\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__39019\,
            I => \N__39014\
        );

    \I__8101\ : InMux
    port map (
            O => \N__39018\,
            I => \N__39011\
        );

    \I__8100\ : InMux
    port map (
            O => \N__39017\,
            I => \N__39008\
        );

    \I__8099\ : Span4Mux_h
    port map (
            O => \N__39014\,
            I => \N__39005\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__39011\,
            I => \N__39002\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__39008\,
            I => \N__38999\
        );

    \I__8096\ : Odrv4
    port map (
            O => \N__39005\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__8095\ : Odrv4
    port map (
            O => \N__39002\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__8094\ : Odrv4
    port map (
            O => \N__38999\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__8093\ : InMux
    port map (
            O => \N__38992\,
            I => \N__38988\
        );

    \I__8092\ : CascadeMux
    port map (
            O => \N__38991\,
            I => \N__38985\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__38988\,
            I => \N__38982\
        );

    \I__8090\ : InMux
    port map (
            O => \N__38985\,
            I => \N__38979\
        );

    \I__8089\ : Span4Mux_v
    port map (
            O => \N__38982\,
            I => \N__38975\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__38979\,
            I => \N__38972\
        );

    \I__8087\ : InMux
    port map (
            O => \N__38978\,
            I => \N__38969\
        );

    \I__8086\ : Odrv4
    port map (
            O => \N__38975\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__8085\ : Odrv4
    port map (
            O => \N__38972\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__38969\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__8083\ : CascadeMux
    port map (
            O => \N__38962\,
            I => \N__38957\
        );

    \I__8082\ : InMux
    port map (
            O => \N__38961\,
            I => \N__38954\
        );

    \I__8081\ : InMux
    port map (
            O => \N__38960\,
            I => \N__38951\
        );

    \I__8080\ : InMux
    port map (
            O => \N__38957\,
            I => \N__38948\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__38954\,
            I => \N__38945\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__38951\,
            I => \N__38940\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__38948\,
            I => \N__38940\
        );

    \I__8076\ : Odrv4
    port map (
            O => \N__38945\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__8075\ : Odrv4
    port map (
            O => \N__38940\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__8074\ : InMux
    port map (
            O => \N__38935\,
            I => \N__38931\
        );

    \I__8073\ : InMux
    port map (
            O => \N__38934\,
            I => \N__38928\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__38931\,
            I => \N__38925\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__38928\,
            I => \N__38922\
        );

    \I__8070\ : Span4Mux_h
    port map (
            O => \N__38925\,
            I => \N__38919\
        );

    \I__8069\ : Span4Mux_h
    port map (
            O => \N__38922\,
            I => \N__38916\
        );

    \I__8068\ : Odrv4
    port map (
            O => \N__38919\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1\
        );

    \I__8067\ : Odrv4
    port map (
            O => \N__38916\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1\
        );

    \I__8066\ : InMux
    port map (
            O => \N__38911\,
            I => \N__38908\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__38908\,
            I => \N__38905\
        );

    \I__8064\ : Span4Mux_h
    port map (
            O => \N__38905\,
            I => \N__38901\
        );

    \I__8063\ : InMux
    port map (
            O => \N__38904\,
            I => \N__38898\
        );

    \I__8062\ : Span4Mux_v
    port map (
            O => \N__38901\,
            I => \N__38894\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__38898\,
            I => \N__38891\
        );

    \I__8060\ : InMux
    port map (
            O => \N__38897\,
            I => \N__38888\
        );

    \I__8059\ : Odrv4
    port map (
            O => \N__38894\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8058\ : Odrv12
    port map (
            O => \N__38891\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__38888\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8056\ : InMux
    port map (
            O => \N__38881\,
            I => \N__38878\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__38878\,
            I => \N__38874\
        );

    \I__8054\ : InMux
    port map (
            O => \N__38877\,
            I => \N__38871\
        );

    \I__8053\ : Span4Mux_v
    port map (
            O => \N__38874\,
            I => \N__38866\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__38871\,
            I => \N__38866\
        );

    \I__8051\ : Odrv4
    port map (
            O => \N__38866\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__8050\ : InMux
    port map (
            O => \N__38863\,
            I => \N__38860\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__38860\,
            I => \N__38856\
        );

    \I__8048\ : InMux
    port map (
            O => \N__38859\,
            I => \N__38853\
        );

    \I__8047\ : Span4Mux_v
    port map (
            O => \N__38856\,
            I => \N__38849\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__38853\,
            I => \N__38846\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38852\,
            I => \N__38843\
        );

    \I__8044\ : Odrv4
    port map (
            O => \N__38849\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8043\ : Odrv12
    port map (
            O => \N__38846\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__38843\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8041\ : InMux
    port map (
            O => \N__38836\,
            I => \N__38833\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__38833\,
            I => \N__38828\
        );

    \I__8039\ : InMux
    port map (
            O => \N__38832\,
            I => \N__38825\
        );

    \I__8038\ : InMux
    port map (
            O => \N__38831\,
            I => \N__38822\
        );

    \I__8037\ : Span4Mux_v
    port map (
            O => \N__38828\,
            I => \N__38817\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__38825\,
            I => \N__38817\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__38822\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__8034\ : Odrv4
    port map (
            O => \N__38817\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__8033\ : CEMux
    port map (
            O => \N__38812\,
            I => \N__38797\
        );

    \I__8032\ : CEMux
    port map (
            O => \N__38811\,
            I => \N__38797\
        );

    \I__8031\ : CEMux
    port map (
            O => \N__38810\,
            I => \N__38797\
        );

    \I__8030\ : CEMux
    port map (
            O => \N__38809\,
            I => \N__38797\
        );

    \I__8029\ : CEMux
    port map (
            O => \N__38808\,
            I => \N__38797\
        );

    \I__8028\ : GlobalMux
    port map (
            O => \N__38797\,
            I => \N__38794\
        );

    \I__8027\ : gio2CtrlBuf
    port map (
            O => \N__38794\,
            I => \delay_measurement_inst.delay_hc_timer.N_302_i_g\
        );

    \I__8026\ : CascadeMux
    port map (
            O => \N__38791\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3_cascade_\
        );

    \I__8025\ : InMux
    port map (
            O => \N__38788\,
            I => \N__38785\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__38785\,
            I => \N__38782\
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__38782\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4\
        );

    \I__8022\ : InMux
    port map (
            O => \N__38779\,
            I => \N__38773\
        );

    \I__8021\ : InMux
    port map (
            O => \N__38778\,
            I => \N__38770\
        );

    \I__8020\ : InMux
    port map (
            O => \N__38777\,
            I => \N__38767\
        );

    \I__8019\ : InMux
    port map (
            O => \N__38776\,
            I => \N__38764\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__38773\,
            I => \N__38757\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__38770\,
            I => \N__38757\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__38767\,
            I => \N__38757\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__38764\,
            I => \N__38754\
        );

    \I__8014\ : Span4Mux_v
    port map (
            O => \N__38757\,
            I => \N__38751\
        );

    \I__8013\ : Span4Mux_h
    port map (
            O => \N__38754\,
            I => \N__38748\
        );

    \I__8012\ : Span4Mux_h
    port map (
            O => \N__38751\,
            I => \N__38745\
        );

    \I__8011\ : Span4Mux_v
    port map (
            O => \N__38748\,
            I => \N__38742\
        );

    \I__8010\ : Odrv4
    port map (
            O => \N__38745\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1\
        );

    \I__8009\ : Odrv4
    port map (
            O => \N__38742\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1\
        );

    \I__8008\ : InMux
    port map (
            O => \N__38737\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__8007\ : InMux
    port map (
            O => \N__38734\,
            I => \N__38731\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__38731\,
            I => \N__38728\
        );

    \I__8005\ : Span4Mux_h
    port map (
            O => \N__38728\,
            I => \N__38725\
        );

    \I__8004\ : Span4Mux_v
    port map (
            O => \N__38725\,
            I => \N__38722\
        );

    \I__8003\ : Odrv4
    port map (
            O => \N__38722\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__8002\ : InMux
    port map (
            O => \N__38719\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__8001\ : InMux
    port map (
            O => \N__38716\,
            I => \N__38713\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__38713\,
            I => \N__38710\
        );

    \I__7999\ : Span4Mux_h
    port map (
            O => \N__38710\,
            I => \N__38707\
        );

    \I__7998\ : Odrv4
    port map (
            O => \N__38707\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__7997\ : InMux
    port map (
            O => \N__38704\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__7996\ : InMux
    port map (
            O => \N__38701\,
            I => \N__38698\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__38698\,
            I => \N__38695\
        );

    \I__7994\ : Span4Mux_h
    port map (
            O => \N__38695\,
            I => \N__38692\
        );

    \I__7993\ : Span4Mux_v
    port map (
            O => \N__38692\,
            I => \N__38689\
        );

    \I__7992\ : Odrv4
    port map (
            O => \N__38689\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__7991\ : InMux
    port map (
            O => \N__38686\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__7990\ : InMux
    port map (
            O => \N__38683\,
            I => \N__38680\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__38680\,
            I => \N__38677\
        );

    \I__7988\ : Span4Mux_h
    port map (
            O => \N__38677\,
            I => \N__38674\
        );

    \I__7987\ : Odrv4
    port map (
            O => \N__38674\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__7986\ : InMux
    port map (
            O => \N__38671\,
            I => \bfn_15_22_0_\
        );

    \I__7985\ : InMux
    port map (
            O => \N__38668\,
            I => \N__38665\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__38665\,
            I => \N__38662\
        );

    \I__7983\ : Odrv4
    port map (
            O => \N__38662\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__7982\ : InMux
    port map (
            O => \N__38659\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__7981\ : InMux
    port map (
            O => \N__38656\,
            I => \N__38653\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__38653\,
            I => \N__38650\
        );

    \I__7979\ : Odrv4
    port map (
            O => \N__38650\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__7978\ : InMux
    port map (
            O => \N__38647\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__7977\ : CascadeMux
    port map (
            O => \N__38644\,
            I => \N__38641\
        );

    \I__7976\ : InMux
    port map (
            O => \N__38641\,
            I => \N__38638\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__38638\,
            I => \N__38635\
        );

    \I__7974\ : Odrv4
    port map (
            O => \N__38635\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__7973\ : InMux
    port map (
            O => \N__38632\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__7972\ : InMux
    port map (
            O => \N__38629\,
            I => \N__38626\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__38626\,
            I => \N__38623\
        );

    \I__7970\ : Span4Mux_h
    port map (
            O => \N__38623\,
            I => \N__38620\
        );

    \I__7969\ : Odrv4
    port map (
            O => \N__38620\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__7968\ : InMux
    port map (
            O => \N__38617\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__7967\ : InMux
    port map (
            O => \N__38614\,
            I => \N__38611\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__38611\,
            I => \N__38608\
        );

    \I__7965\ : Span4Mux_h
    port map (
            O => \N__38608\,
            I => \N__38605\
        );

    \I__7964\ : Span4Mux_v
    port map (
            O => \N__38605\,
            I => \N__38602\
        );

    \I__7963\ : Odrv4
    port map (
            O => \N__38602\,
            I => \current_shift_inst.un38_control_input_0_s1_12\
        );

    \I__7962\ : InMux
    port map (
            O => \N__38599\,
            I => \current_shift_inst.un38_control_input_cry_11_s1\
        );

    \I__7961\ : InMux
    port map (
            O => \N__38596\,
            I => \current_shift_inst.un38_control_input_cry_12_s1\
        );

    \I__7960\ : InMux
    port map (
            O => \N__38593\,
            I => \N__38590\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__38590\,
            I => \N__38587\
        );

    \I__7958\ : Span4Mux_h
    port map (
            O => \N__38587\,
            I => \N__38584\
        );

    \I__7957\ : Span4Mux_v
    port map (
            O => \N__38584\,
            I => \N__38581\
        );

    \I__7956\ : Odrv4
    port map (
            O => \N__38581\,
            I => \current_shift_inst.un38_control_input_0_s1_14\
        );

    \I__7955\ : InMux
    port map (
            O => \N__38578\,
            I => \current_shift_inst.un38_control_input_cry_13_s1\
        );

    \I__7954\ : InMux
    port map (
            O => \N__38575\,
            I => \N__38572\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__38572\,
            I => \N__38569\
        );

    \I__7952\ : Span4Mux_h
    port map (
            O => \N__38569\,
            I => \N__38566\
        );

    \I__7951\ : Span4Mux_v
    port map (
            O => \N__38566\,
            I => \N__38563\
        );

    \I__7950\ : Odrv4
    port map (
            O => \N__38563\,
            I => \current_shift_inst.un38_control_input_0_s1_15\
        );

    \I__7949\ : InMux
    port map (
            O => \N__38560\,
            I => \current_shift_inst.un38_control_input_cry_14_s1\
        );

    \I__7948\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38554\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__38554\,
            I => \N__38551\
        );

    \I__7946\ : Span4Mux_h
    port map (
            O => \N__38551\,
            I => \N__38548\
        );

    \I__7945\ : Span4Mux_v
    port map (
            O => \N__38548\,
            I => \N__38545\
        );

    \I__7944\ : Odrv4
    port map (
            O => \N__38545\,
            I => \current_shift_inst.un38_control_input_0_s1_16\
        );

    \I__7943\ : InMux
    port map (
            O => \N__38542\,
            I => \bfn_15_21_0_\
        );

    \I__7942\ : InMux
    port map (
            O => \N__38539\,
            I => \N__38536\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__38536\,
            I => \N__38533\
        );

    \I__7940\ : Span4Mux_h
    port map (
            O => \N__38533\,
            I => \N__38530\
        );

    \I__7939\ : Span4Mux_v
    port map (
            O => \N__38530\,
            I => \N__38527\
        );

    \I__7938\ : Odrv4
    port map (
            O => \N__38527\,
            I => \current_shift_inst.un38_control_input_0_s1_17\
        );

    \I__7937\ : InMux
    port map (
            O => \N__38524\,
            I => \current_shift_inst.un38_control_input_cry_16_s1\
        );

    \I__7936\ : InMux
    port map (
            O => \N__38521\,
            I => \N__38518\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__38518\,
            I => \N__38515\
        );

    \I__7934\ : Span4Mux_v
    port map (
            O => \N__38515\,
            I => \N__38512\
        );

    \I__7933\ : Span4Mux_v
    port map (
            O => \N__38512\,
            I => \N__38509\
        );

    \I__7932\ : Odrv4
    port map (
            O => \N__38509\,
            I => \current_shift_inst.un38_control_input_0_s1_18\
        );

    \I__7931\ : InMux
    port map (
            O => \N__38506\,
            I => \current_shift_inst.un38_control_input_cry_17_s1\
        );

    \I__7930\ : InMux
    port map (
            O => \N__38503\,
            I => \N__38500\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__38500\,
            I => \N__38497\
        );

    \I__7928\ : Span4Mux_h
    port map (
            O => \N__38497\,
            I => \N__38494\
        );

    \I__7927\ : Span4Mux_v
    port map (
            O => \N__38494\,
            I => \N__38491\
        );

    \I__7926\ : Odrv4
    port map (
            O => \N__38491\,
            I => \current_shift_inst.un38_control_input_0_s1_19\
        );

    \I__7925\ : InMux
    port map (
            O => \N__38488\,
            I => \current_shift_inst.un38_control_input_cry_18_s1\
        );

    \I__7924\ : InMux
    port map (
            O => \N__38485\,
            I => \N__38482\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__38482\,
            I => \N__38479\
        );

    \I__7922\ : Span4Mux_h
    port map (
            O => \N__38479\,
            I => \N__38476\
        );

    \I__7921\ : Span4Mux_v
    port map (
            O => \N__38476\,
            I => \N__38473\
        );

    \I__7920\ : Odrv4
    port map (
            O => \N__38473\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__7919\ : InMux
    port map (
            O => \N__38470\,
            I => \N__38467\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__38467\,
            I => \current_shift_inst.un38_control_input_0_s1_6\
        );

    \I__7917\ : InMux
    port map (
            O => \N__38464\,
            I => \current_shift_inst.un38_control_input_cry_5_s1\
        );

    \I__7916\ : InMux
    port map (
            O => \N__38461\,
            I => \N__38458\
        );

    \I__7915\ : LocalMux
    port map (
            O => \N__38458\,
            I => \N__38455\
        );

    \I__7914\ : Odrv4
    port map (
            O => \N__38455\,
            I => \current_shift_inst.un38_control_input_0_s1_7\
        );

    \I__7913\ : InMux
    port map (
            O => \N__38452\,
            I => \current_shift_inst.un38_control_input_cry_6_s1\
        );

    \I__7912\ : InMux
    port map (
            O => \N__38449\,
            I => \N__38446\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__38446\,
            I => \N__38443\
        );

    \I__7910\ : Span4Mux_h
    port map (
            O => \N__38443\,
            I => \N__38440\
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__38440\,
            I => \current_shift_inst.un38_control_input_0_s1_8\
        );

    \I__7908\ : InMux
    port map (
            O => \N__38437\,
            I => \bfn_15_20_0_\
        );

    \I__7907\ : InMux
    port map (
            O => \N__38434\,
            I => \N__38431\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__38431\,
            I => \N__38428\
        );

    \I__7905\ : Span4Mux_h
    port map (
            O => \N__38428\,
            I => \N__38425\
        );

    \I__7904\ : Odrv4
    port map (
            O => \N__38425\,
            I => \current_shift_inst.un38_control_input_0_s1_9\
        );

    \I__7903\ : InMux
    port map (
            O => \N__38422\,
            I => \current_shift_inst.un38_control_input_cry_8_s1\
        );

    \I__7902\ : InMux
    port map (
            O => \N__38419\,
            I => \N__38416\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__38416\,
            I => \N__38413\
        );

    \I__7900\ : Span4Mux_h
    port map (
            O => \N__38413\,
            I => \N__38410\
        );

    \I__7899\ : Span4Mux_v
    port map (
            O => \N__38410\,
            I => \N__38407\
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__38407\,
            I => \current_shift_inst.un38_control_input_0_s1_10\
        );

    \I__7897\ : InMux
    port map (
            O => \N__38404\,
            I => \current_shift_inst.un38_control_input_cry_9_s1\
        );

    \I__7896\ : InMux
    port map (
            O => \N__38401\,
            I => \current_shift_inst.un38_control_input_cry_10_s1\
        );

    \I__7895\ : InMux
    port map (
            O => \N__38398\,
            I => \N__38395\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__38395\,
            I => \N__38369\
        );

    \I__7893\ : InMux
    port map (
            O => \N__38394\,
            I => \N__38355\
        );

    \I__7892\ : InMux
    port map (
            O => \N__38393\,
            I => \N__38355\
        );

    \I__7891\ : InMux
    port map (
            O => \N__38392\,
            I => \N__38355\
        );

    \I__7890\ : InMux
    port map (
            O => \N__38391\,
            I => \N__38346\
        );

    \I__7889\ : InMux
    port map (
            O => \N__38390\,
            I => \N__38346\
        );

    \I__7888\ : InMux
    port map (
            O => \N__38389\,
            I => \N__38346\
        );

    \I__7887\ : InMux
    port map (
            O => \N__38388\,
            I => \N__38346\
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__38387\,
            I => \N__38343\
        );

    \I__7885\ : CascadeMux
    port map (
            O => \N__38386\,
            I => \N__38340\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__38385\,
            I => \N__38336\
        );

    \I__7883\ : CascadeMux
    port map (
            O => \N__38384\,
            I => \N__38333\
        );

    \I__7882\ : CascadeMux
    port map (
            O => \N__38383\,
            I => \N__38330\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__38382\,
            I => \N__38327\
        );

    \I__7880\ : CascadeMux
    port map (
            O => \N__38381\,
            I => \N__38323\
        );

    \I__7879\ : CascadeMux
    port map (
            O => \N__38380\,
            I => \N__38320\
        );

    \I__7878\ : CascadeMux
    port map (
            O => \N__38379\,
            I => \N__38317\
        );

    \I__7877\ : CascadeMux
    port map (
            O => \N__38378\,
            I => \N__38314\
        );

    \I__7876\ : CascadeMux
    port map (
            O => \N__38377\,
            I => \N__38311\
        );

    \I__7875\ : CascadeMux
    port map (
            O => \N__38376\,
            I => \N__38308\
        );

    \I__7874\ : CascadeMux
    port map (
            O => \N__38375\,
            I => \N__38305\
        );

    \I__7873\ : CascadeMux
    port map (
            O => \N__38374\,
            I => \N__38302\
        );

    \I__7872\ : CascadeMux
    port map (
            O => \N__38373\,
            I => \N__38299\
        );

    \I__7871\ : CascadeMux
    port map (
            O => \N__38372\,
            I => \N__38296\
        );

    \I__7870\ : Span4Mux_s2_h
    port map (
            O => \N__38369\,
            I => \N__38276\
        );

    \I__7869\ : InMux
    port map (
            O => \N__38368\,
            I => \N__38269\
        );

    \I__7868\ : InMux
    port map (
            O => \N__38367\,
            I => \N__38269\
        );

    \I__7867\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38269\
        );

    \I__7866\ : InMux
    port map (
            O => \N__38365\,
            I => \N__38260\
        );

    \I__7865\ : InMux
    port map (
            O => \N__38364\,
            I => \N__38260\
        );

    \I__7864\ : InMux
    port map (
            O => \N__38363\,
            I => \N__38260\
        );

    \I__7863\ : InMux
    port map (
            O => \N__38362\,
            I => \N__38260\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__38355\,
            I => \N__38255\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__38346\,
            I => \N__38255\
        );

    \I__7860\ : InMux
    port map (
            O => \N__38343\,
            I => \N__38252\
        );

    \I__7859\ : InMux
    port map (
            O => \N__38340\,
            I => \N__38247\
        );

    \I__7858\ : InMux
    port map (
            O => \N__38339\,
            I => \N__38247\
        );

    \I__7857\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38242\
        );

    \I__7856\ : InMux
    port map (
            O => \N__38333\,
            I => \N__38242\
        );

    \I__7855\ : InMux
    port map (
            O => \N__38330\,
            I => \N__38231\
        );

    \I__7854\ : InMux
    port map (
            O => \N__38327\,
            I => \N__38231\
        );

    \I__7853\ : InMux
    port map (
            O => \N__38326\,
            I => \N__38231\
        );

    \I__7852\ : InMux
    port map (
            O => \N__38323\,
            I => \N__38231\
        );

    \I__7851\ : InMux
    port map (
            O => \N__38320\,
            I => \N__38231\
        );

    \I__7850\ : InMux
    port map (
            O => \N__38317\,
            I => \N__38222\
        );

    \I__7849\ : InMux
    port map (
            O => \N__38314\,
            I => \N__38222\
        );

    \I__7848\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38222\
        );

    \I__7847\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38222\
        );

    \I__7846\ : InMux
    port map (
            O => \N__38305\,
            I => \N__38213\
        );

    \I__7845\ : InMux
    port map (
            O => \N__38302\,
            I => \N__38213\
        );

    \I__7844\ : InMux
    port map (
            O => \N__38299\,
            I => \N__38213\
        );

    \I__7843\ : InMux
    port map (
            O => \N__38296\,
            I => \N__38213\
        );

    \I__7842\ : CascadeMux
    port map (
            O => \N__38295\,
            I => \N__38210\
        );

    \I__7841\ : CascadeMux
    port map (
            O => \N__38294\,
            I => \N__38207\
        );

    \I__7840\ : CascadeMux
    port map (
            O => \N__38293\,
            I => \N__38204\
        );

    \I__7839\ : CascadeMux
    port map (
            O => \N__38292\,
            I => \N__38201\
        );

    \I__7838\ : CascadeMux
    port map (
            O => \N__38291\,
            I => \N__38197\
        );

    \I__7837\ : CascadeMux
    port map (
            O => \N__38290\,
            I => \N__38194\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__38289\,
            I => \N__38191\
        );

    \I__7835\ : InMux
    port map (
            O => \N__38288\,
            I => \N__38188\
        );

    \I__7834\ : InMux
    port map (
            O => \N__38287\,
            I => \N__38185\
        );

    \I__7833\ : CascadeMux
    port map (
            O => \N__38286\,
            I => \N__38182\
        );

    \I__7832\ : CascadeMux
    port map (
            O => \N__38285\,
            I => \N__38179\
        );

    \I__7831\ : CascadeMux
    port map (
            O => \N__38284\,
            I => \N__38176\
        );

    \I__7830\ : CascadeMux
    port map (
            O => \N__38283\,
            I => \N__38173\
        );

    \I__7829\ : CascadeMux
    port map (
            O => \N__38282\,
            I => \N__38170\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__38281\,
            I => \N__38167\
        );

    \I__7827\ : CascadeMux
    port map (
            O => \N__38280\,
            I => \N__38164\
        );

    \I__7826\ : InMux
    port map (
            O => \N__38279\,
            I => \N__38159\
        );

    \I__7825\ : Span4Mux_h
    port map (
            O => \N__38276\,
            I => \N__38156\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__38269\,
            I => \N__38151\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__38260\,
            I => \N__38151\
        );

    \I__7822\ : Span4Mux_s3_h
    port map (
            O => \N__38255\,
            I => \N__38148\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__38252\,
            I => \N__38143\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__38247\,
            I => \N__38143\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__38242\,
            I => \N__38134\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__38231\,
            I => \N__38134\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__38222\,
            I => \N__38134\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__38213\,
            I => \N__38134\
        );

    \I__7815\ : InMux
    port map (
            O => \N__38210\,
            I => \N__38127\
        );

    \I__7814\ : InMux
    port map (
            O => \N__38207\,
            I => \N__38127\
        );

    \I__7813\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38127\
        );

    \I__7812\ : InMux
    port map (
            O => \N__38201\,
            I => \N__38116\
        );

    \I__7811\ : InMux
    port map (
            O => \N__38200\,
            I => \N__38116\
        );

    \I__7810\ : InMux
    port map (
            O => \N__38197\,
            I => \N__38116\
        );

    \I__7809\ : InMux
    port map (
            O => \N__38194\,
            I => \N__38116\
        );

    \I__7808\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38116\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__38188\,
            I => \N__38113\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__38185\,
            I => \N__38110\
        );

    \I__7805\ : InMux
    port map (
            O => \N__38182\,
            I => \N__38103\
        );

    \I__7804\ : InMux
    port map (
            O => \N__38179\,
            I => \N__38103\
        );

    \I__7803\ : InMux
    port map (
            O => \N__38176\,
            I => \N__38103\
        );

    \I__7802\ : InMux
    port map (
            O => \N__38173\,
            I => \N__38094\
        );

    \I__7801\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38094\
        );

    \I__7800\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38094\
        );

    \I__7799\ : InMux
    port map (
            O => \N__38164\,
            I => \N__38094\
        );

    \I__7798\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38091\
        );

    \I__7797\ : InMux
    port map (
            O => \N__38162\,
            I => \N__38088\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__38159\,
            I => \N__38083\
        );

    \I__7795\ : Span4Mux_v
    port map (
            O => \N__38156\,
            I => \N__38078\
        );

    \I__7794\ : Span4Mux_s2_h
    port map (
            O => \N__38151\,
            I => \N__38078\
        );

    \I__7793\ : Span4Mux_v
    port map (
            O => \N__38148\,
            I => \N__38073\
        );

    \I__7792\ : Span4Mux_s3_h
    port map (
            O => \N__38143\,
            I => \N__38073\
        );

    \I__7791\ : Span4Mux_v
    port map (
            O => \N__38134\,
            I => \N__38070\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__38127\,
            I => \N__38065\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__38116\,
            I => \N__38065\
        );

    \I__7788\ : Span4Mux_v
    port map (
            O => \N__38113\,
            I => \N__38060\
        );

    \I__7787\ : Span4Mux_v
    port map (
            O => \N__38110\,
            I => \N__38060\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__38103\,
            I => \N__38055\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__38094\,
            I => \N__38055\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__38091\,
            I => \N__38052\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__38088\,
            I => \N__38049\
        );

    \I__7782\ : InMux
    port map (
            O => \N__38087\,
            I => \N__38046\
        );

    \I__7781\ : InMux
    port map (
            O => \N__38086\,
            I => \N__38043\
        );

    \I__7780\ : Span12Mux_s2_h
    port map (
            O => \N__38083\,
            I => \N__38038\
        );

    \I__7779\ : Sp12to4
    port map (
            O => \N__38078\,
            I => \N__38038\
        );

    \I__7778\ : Sp12to4
    port map (
            O => \N__38073\,
            I => \N__38035\
        );

    \I__7777\ : Sp12to4
    port map (
            O => \N__38070\,
            I => \N__38028\
        );

    \I__7776\ : Span12Mux_s10_h
    port map (
            O => \N__38065\,
            I => \N__38028\
        );

    \I__7775\ : Sp12to4
    port map (
            O => \N__38060\,
            I => \N__38028\
        );

    \I__7774\ : Span12Mux_v
    port map (
            O => \N__38055\,
            I => \N__38023\
        );

    \I__7773\ : Span12Mux_s10_h
    port map (
            O => \N__38052\,
            I => \N__38023\
        );

    \I__7772\ : Span4Mux_s3_h
    port map (
            O => \N__38049\,
            I => \N__38020\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__38046\,
            I => \N__38015\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__38043\,
            I => \N__38015\
        );

    \I__7769\ : Span12Mux_v
    port map (
            O => \N__38038\,
            I => \N__38012\
        );

    \I__7768\ : Span12Mux_v
    port map (
            O => \N__38035\,
            I => \N__38001\
        );

    \I__7767\ : Span12Mux_h
    port map (
            O => \N__38028\,
            I => \N__38001\
        );

    \I__7766\ : Span12Mux_h
    port map (
            O => \N__38023\,
            I => \N__38001\
        );

    \I__7765\ : Sp12to4
    port map (
            O => \N__38020\,
            I => \N__38001\
        );

    \I__7764\ : Span12Mux_s3_h
    port map (
            O => \N__38015\,
            I => \N__38001\
        );

    \I__7763\ : Odrv12
    port map (
            O => \N__38012\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7762\ : Odrv12
    port map (
            O => \N__38001\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7761\ : InMux
    port map (
            O => \N__37996\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__7760\ : InMux
    port map (
            O => \N__37993\,
            I => \N__37989\
        );

    \I__7759\ : InMux
    port map (
            O => \N__37992\,
            I => \N__37986\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__37989\,
            I => \N__37983\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__37986\,
            I => \N__37978\
        );

    \I__7756\ : Span4Mux_h
    port map (
            O => \N__37983\,
            I => \N__37978\
        );

    \I__7755\ : Odrv4
    port map (
            O => \N__37978\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__7754\ : CascadeMux
    port map (
            O => \N__37975\,
            I => \N__37971\
        );

    \I__7753\ : CascadeMux
    port map (
            O => \N__37974\,
            I => \N__37968\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37971\,
            I => \N__37965\
        );

    \I__7751\ : InMux
    port map (
            O => \N__37968\,
            I => \N__37962\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__37965\,
            I => \N__37959\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__37962\,
            I => \N__37956\
        );

    \I__7748\ : Odrv4
    port map (
            O => \N__37959\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__7747\ : Odrv12
    port map (
            O => \N__37956\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__7746\ : InMux
    port map (
            O => \N__37951\,
            I => \N__37948\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__37948\,
            I => \N__37945\
        );

    \I__7744\ : Span4Mux_h
    port map (
            O => \N__37945\,
            I => \N__37942\
        );

    \I__7743\ : Odrv4
    port map (
            O => \N__37942\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__7742\ : InMux
    port map (
            O => \N__37939\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__7741\ : CascadeMux
    port map (
            O => \N__37936\,
            I => \N__37928\
        );

    \I__7740\ : CascadeMux
    port map (
            O => \N__37935\,
            I => \N__37923\
        );

    \I__7739\ : InMux
    port map (
            O => \N__37934\,
            I => \N__37916\
        );

    \I__7738\ : InMux
    port map (
            O => \N__37933\,
            I => \N__37916\
        );

    \I__7737\ : InMux
    port map (
            O => \N__37932\,
            I => \N__37916\
        );

    \I__7736\ : CascadeMux
    port map (
            O => \N__37931\,
            I => \N__37913\
        );

    \I__7735\ : InMux
    port map (
            O => \N__37928\,
            I => \N__37905\
        );

    \I__7734\ : InMux
    port map (
            O => \N__37927\,
            I => \N__37900\
        );

    \I__7733\ : InMux
    port map (
            O => \N__37926\,
            I => \N__37900\
        );

    \I__7732\ : InMux
    port map (
            O => \N__37923\,
            I => \N__37897\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__37916\,
            I => \N__37894\
        );

    \I__7730\ : InMux
    port map (
            O => \N__37913\,
            I => \N__37881\
        );

    \I__7729\ : InMux
    port map (
            O => \N__37912\,
            I => \N__37881\
        );

    \I__7728\ : InMux
    port map (
            O => \N__37911\,
            I => \N__37881\
        );

    \I__7727\ : InMux
    port map (
            O => \N__37910\,
            I => \N__37881\
        );

    \I__7726\ : InMux
    port map (
            O => \N__37909\,
            I => \N__37881\
        );

    \I__7725\ : InMux
    port map (
            O => \N__37908\,
            I => \N__37881\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__37905\,
            I => \N__37878\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__37900\,
            I => \N__37873\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__37897\,
            I => \N__37873\
        );

    \I__7721\ : Span4Mux_h
    port map (
            O => \N__37894\,
            I => \N__37870\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__37881\,
            I => \N__37867\
        );

    \I__7719\ : Span4Mux_h
    port map (
            O => \N__37878\,
            I => \N__37864\
        );

    \I__7718\ : Span4Mux_h
    port map (
            O => \N__37873\,
            I => \N__37861\
        );

    \I__7717\ : Odrv4
    port map (
            O => \N__37870\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__7716\ : Odrv12
    port map (
            O => \N__37867\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__7715\ : Odrv4
    port map (
            O => \N__37864\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__7714\ : Odrv4
    port map (
            O => \N__37861\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__7713\ : CascadeMux
    port map (
            O => \N__37852\,
            I => \N__37849\
        );

    \I__7712\ : InMux
    port map (
            O => \N__37849\,
            I => \N__37846\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__37846\,
            I => \N__37840\
        );

    \I__7710\ : InMux
    port map (
            O => \N__37845\,
            I => \N__37837\
        );

    \I__7709\ : InMux
    port map (
            O => \N__37844\,
            I => \N__37832\
        );

    \I__7708\ : InMux
    port map (
            O => \N__37843\,
            I => \N__37832\
        );

    \I__7707\ : Span4Mux_h
    port map (
            O => \N__37840\,
            I => \N__37827\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__37837\,
            I => \N__37827\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__37832\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__7704\ : Odrv4
    port map (
            O => \N__37827\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__7703\ : InMux
    port map (
            O => \N__37822\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__7702\ : InMux
    port map (
            O => \N__37819\,
            I => \N__37816\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__37816\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__7700\ : InMux
    port map (
            O => \N__37813\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__7699\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37807\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__37807\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__7697\ : InMux
    port map (
            O => \N__37804\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__7696\ : InMux
    port map (
            O => \N__37801\,
            I => \N__37798\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__37798\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__7694\ : InMux
    port map (
            O => \N__37795\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__7693\ : CascadeMux
    port map (
            O => \N__37792\,
            I => \N__37789\
        );

    \I__7692\ : InMux
    port map (
            O => \N__37789\,
            I => \N__37786\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__37786\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__7690\ : InMux
    port map (
            O => \N__37783\,
            I => \bfn_15_14_0_\
        );

    \I__7689\ : InMux
    port map (
            O => \N__37780\,
            I => \N__37777\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__37777\,
            I => \N__37774\
        );

    \I__7687\ : Odrv12
    port map (
            O => \N__37774\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__7686\ : InMux
    port map (
            O => \N__37771\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__7685\ : InMux
    port map (
            O => \N__37768\,
            I => \N__37765\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__37765\,
            I => \N__37762\
        );

    \I__7683\ : Odrv4
    port map (
            O => \N__37762\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__7682\ : InMux
    port map (
            O => \N__37759\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__7681\ : CascadeMux
    port map (
            O => \N__37756\,
            I => \N__37753\
        );

    \I__7680\ : InMux
    port map (
            O => \N__37753\,
            I => \N__37750\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__37750\,
            I => \N__37747\
        );

    \I__7678\ : Span4Mux_v
    port map (
            O => \N__37747\,
            I => \N__37744\
        );

    \I__7677\ : Odrv4
    port map (
            O => \N__37744\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\
        );

    \I__7676\ : InMux
    port map (
            O => \N__37741\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__7675\ : InMux
    port map (
            O => \N__37738\,
            I => \N__37733\
        );

    \I__7674\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37728\
        );

    \I__7673\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37725\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__37733\,
            I => \N__37722\
        );

    \I__7671\ : InMux
    port map (
            O => \N__37732\,
            I => \N__37717\
        );

    \I__7670\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37717\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__37728\,
            I => \N__37712\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__37725\,
            I => \N__37712\
        );

    \I__7667\ : Span4Mux_v
    port map (
            O => \N__37722\,
            I => \N__37705\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__37717\,
            I => \N__37705\
        );

    \I__7665\ : Span4Mux_v
    port map (
            O => \N__37712\,
            I => \N__37705\
        );

    \I__7664\ : Odrv4
    port map (
            O => \N__37705\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__7663\ : InMux
    port map (
            O => \N__37702\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__7662\ : CascadeMux
    port map (
            O => \N__37699\,
            I => \N__37696\
        );

    \I__7661\ : InMux
    port map (
            O => \N__37696\,
            I => \N__37687\
        );

    \I__7660\ : InMux
    port map (
            O => \N__37695\,
            I => \N__37687\
        );

    \I__7659\ : CascadeMux
    port map (
            O => \N__37694\,
            I => \N__37683\
        );

    \I__7658\ : InMux
    port map (
            O => \N__37693\,
            I => \N__37680\
        );

    \I__7657\ : InMux
    port map (
            O => \N__37692\,
            I => \N__37677\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__37687\,
            I => \N__37674\
        );

    \I__7655\ : InMux
    port map (
            O => \N__37686\,
            I => \N__37669\
        );

    \I__7654\ : InMux
    port map (
            O => \N__37683\,
            I => \N__37669\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__37680\,
            I => \N__37660\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__37677\,
            I => \N__37660\
        );

    \I__7651\ : Span4Mux_v
    port map (
            O => \N__37674\,
            I => \N__37660\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__37669\,
            I => \N__37660\
        );

    \I__7649\ : Span4Mux_v
    port map (
            O => \N__37660\,
            I => \N__37657\
        );

    \I__7648\ : Odrv4
    port map (
            O => \N__37657\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__7647\ : InMux
    port map (
            O => \N__37654\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__7646\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37648\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__37648\,
            I => \N__37643\
        );

    \I__7644\ : InMux
    port map (
            O => \N__37647\,
            I => \N__37640\
        );

    \I__7643\ : InMux
    port map (
            O => \N__37646\,
            I => \N__37637\
        );

    \I__7642\ : Span4Mux_v
    port map (
            O => \N__37643\,
            I => \N__37634\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__37640\,
            I => \N__37629\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__37637\,
            I => \N__37629\
        );

    \I__7639\ : Span4Mux_h
    port map (
            O => \N__37634\,
            I => \N__37626\
        );

    \I__7638\ : Span4Mux_v
    port map (
            O => \N__37629\,
            I => \N__37623\
        );

    \I__7637\ : Odrv4
    port map (
            O => \N__37626\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__7636\ : Odrv4
    port map (
            O => \N__37623\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__7635\ : InMux
    port map (
            O => \N__37618\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__7634\ : CascadeMux
    port map (
            O => \N__37615\,
            I => \N__37611\
        );

    \I__7633\ : InMux
    port map (
            O => \N__37614\,
            I => \N__37607\
        );

    \I__7632\ : InMux
    port map (
            O => \N__37611\,
            I => \N__37604\
        );

    \I__7631\ : InMux
    port map (
            O => \N__37610\,
            I => \N__37601\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__37607\,
            I => \N__37598\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__37604\,
            I => \N__37595\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__37601\,
            I => \N__37592\
        );

    \I__7627\ : Span4Mux_v
    port map (
            O => \N__37598\,
            I => \N__37589\
        );

    \I__7626\ : Span4Mux_h
    port map (
            O => \N__37595\,
            I => \N__37586\
        );

    \I__7625\ : Span4Mux_h
    port map (
            O => \N__37592\,
            I => \N__37583\
        );

    \I__7624\ : Odrv4
    port map (
            O => \N__37589\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__7623\ : Odrv4
    port map (
            O => \N__37586\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__7622\ : Odrv4
    port map (
            O => \N__37583\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__7621\ : InMux
    port map (
            O => \N__37576\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__7620\ : InMux
    port map (
            O => \N__37573\,
            I => \N__37568\
        );

    \I__7619\ : InMux
    port map (
            O => \N__37572\,
            I => \N__37565\
        );

    \I__7618\ : InMux
    port map (
            O => \N__37571\,
            I => \N__37562\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__37568\,
            I => \N__37559\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__37565\,
            I => \N__37556\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__37562\,
            I => \N__37553\
        );

    \I__7614\ : Span4Mux_v
    port map (
            O => \N__37559\,
            I => \N__37550\
        );

    \I__7613\ : Span4Mux_h
    port map (
            O => \N__37556\,
            I => \N__37547\
        );

    \I__7612\ : Span4Mux_h
    port map (
            O => \N__37553\,
            I => \N__37544\
        );

    \I__7611\ : Odrv4
    port map (
            O => \N__37550\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__7610\ : Odrv4
    port map (
            O => \N__37547\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__7609\ : Odrv4
    port map (
            O => \N__37544\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__7608\ : InMux
    port map (
            O => \N__37537\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__7607\ : InMux
    port map (
            O => \N__37534\,
            I => \N__37529\
        );

    \I__7606\ : InMux
    port map (
            O => \N__37533\,
            I => \N__37526\
        );

    \I__7605\ : CascadeMux
    port map (
            O => \N__37532\,
            I => \N__37523\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__37529\,
            I => \N__37520\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__37526\,
            I => \N__37517\
        );

    \I__7602\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37514\
        );

    \I__7601\ : Span4Mux_v
    port map (
            O => \N__37520\,
            I => \N__37511\
        );

    \I__7600\ : Span4Mux_h
    port map (
            O => \N__37517\,
            I => \N__37508\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__37514\,
            I => \N__37505\
        );

    \I__7598\ : Odrv4
    port map (
            O => \N__37511\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__7597\ : Odrv4
    port map (
            O => \N__37508\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__7596\ : Odrv12
    port map (
            O => \N__37505\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__7595\ : InMux
    port map (
            O => \N__37498\,
            I => \bfn_15_13_0_\
        );

    \I__7594\ : InMux
    port map (
            O => \N__37495\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__7593\ : InMux
    port map (
            O => \N__37492\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__7592\ : InMux
    port map (
            O => \N__37489\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__7591\ : InMux
    port map (
            O => \N__37486\,
            I => \N__37475\
        );

    \I__7590\ : InMux
    port map (
            O => \N__37485\,
            I => \N__37475\
        );

    \I__7589\ : InMux
    port map (
            O => \N__37484\,
            I => \N__37465\
        );

    \I__7588\ : InMux
    port map (
            O => \N__37483\,
            I => \N__37465\
        );

    \I__7587\ : InMux
    port map (
            O => \N__37482\,
            I => \N__37465\
        );

    \I__7586\ : InMux
    port map (
            O => \N__37481\,
            I => \N__37465\
        );

    \I__7585\ : InMux
    port map (
            O => \N__37480\,
            I => \N__37462\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__37475\,
            I => \N__37459\
        );

    \I__7583\ : InMux
    port map (
            O => \N__37474\,
            I => \N__37456\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__37465\,
            I => \N__37451\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__37462\,
            I => \N__37451\
        );

    \I__7580\ : Span4Mux_v
    port map (
            O => \N__37459\,
            I => \N__37446\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__37456\,
            I => \N__37446\
        );

    \I__7578\ : Span4Mux_v
    port map (
            O => \N__37451\,
            I => \N__37443\
        );

    \I__7577\ : Span4Mux_h
    port map (
            O => \N__37446\,
            I => \N__37440\
        );

    \I__7576\ : Odrv4
    port map (
            O => \N__37443\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__7575\ : Odrv4
    port map (
            O => \N__37440\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__7574\ : InMux
    port map (
            O => \N__37435\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__7573\ : InMux
    port map (
            O => \N__37432\,
            I => \N__37428\
        );

    \I__7572\ : InMux
    port map (
            O => \N__37431\,
            I => \N__37425\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__37428\,
            I => \N__37422\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__37425\,
            I => \N__37419\
        );

    \I__7569\ : Span4Mux_v
    port map (
            O => \N__37422\,
            I => \N__37416\
        );

    \I__7568\ : Span4Mux_v
    port map (
            O => \N__37419\,
            I => \N__37413\
        );

    \I__7567\ : Odrv4
    port map (
            O => \N__37416\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__7566\ : Odrv4
    port map (
            O => \N__37413\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__7565\ : InMux
    port map (
            O => \N__37408\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__7564\ : InMux
    port map (
            O => \N__37405\,
            I => \N__37401\
        );

    \I__7563\ : InMux
    port map (
            O => \N__37404\,
            I => \N__37398\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__37401\,
            I => \N__37395\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__37398\,
            I => \N__37392\
        );

    \I__7560\ : Span4Mux_v
    port map (
            O => \N__37395\,
            I => \N__37389\
        );

    \I__7559\ : Odrv12
    port map (
            O => \N__37392\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__7558\ : Odrv4
    port map (
            O => \N__37389\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__7557\ : InMux
    port map (
            O => \N__37384\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__37381\,
            I => \N__37377\
        );

    \I__7555\ : InMux
    port map (
            O => \N__37380\,
            I => \N__37372\
        );

    \I__7554\ : InMux
    port map (
            O => \N__37377\,
            I => \N__37372\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__37372\,
            I => \N__37366\
        );

    \I__7552\ : InMux
    port map (
            O => \N__37371\,
            I => \N__37363\
        );

    \I__7551\ : InMux
    port map (
            O => \N__37370\,
            I => \N__37360\
        );

    \I__7550\ : InMux
    port map (
            O => \N__37369\,
            I => \N__37357\
        );

    \I__7549\ : Span4Mux_h
    port map (
            O => \N__37366\,
            I => \N__37354\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__37363\,
            I => \N__37349\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__37360\,
            I => \N__37349\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__37357\,
            I => \N__37346\
        );

    \I__7545\ : Span4Mux_h
    port map (
            O => \N__37354\,
            I => \N__37343\
        );

    \I__7544\ : Span4Mux_h
    port map (
            O => \N__37349\,
            I => \N__37340\
        );

    \I__7543\ : Span4Mux_h
    port map (
            O => \N__37346\,
            I => \N__37337\
        );

    \I__7542\ : Odrv4
    port map (
            O => \N__37343\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__7541\ : Odrv4
    port map (
            O => \N__37340\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__7540\ : Odrv4
    port map (
            O => \N__37337\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__7539\ : InMux
    port map (
            O => \N__37330\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__7538\ : InMux
    port map (
            O => \N__37327\,
            I => \N__37324\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__37324\,
            I => \N__37320\
        );

    \I__7536\ : InMux
    port map (
            O => \N__37323\,
            I => \N__37317\
        );

    \I__7535\ : Span4Mux_v
    port map (
            O => \N__37320\,
            I => \N__37312\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__37317\,
            I => \N__37312\
        );

    \I__7533\ : Span4Mux_h
    port map (
            O => \N__37312\,
            I => \N__37309\
        );

    \I__7532\ : Odrv4
    port map (
            O => \N__37309\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__7531\ : InMux
    port map (
            O => \N__37306\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__7530\ : InMux
    port map (
            O => \N__37303\,
            I => \N__37300\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__37300\,
            I => \N__37296\
        );

    \I__7528\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37293\
        );

    \I__7527\ : Span12Mux_v
    port map (
            O => \N__37296\,
            I => \N__37288\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__37293\,
            I => \N__37288\
        );

    \I__7525\ : Odrv12
    port map (
            O => \N__37288\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__7524\ : InMux
    port map (
            O => \N__37285\,
            I => \bfn_15_12_0_\
        );

    \I__7523\ : InMux
    port map (
            O => \N__37282\,
            I => \N__37279\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__37279\,
            I => \N__37275\
        );

    \I__7521\ : InMux
    port map (
            O => \N__37278\,
            I => \N__37272\
        );

    \I__7520\ : Span4Mux_h
    port map (
            O => \N__37275\,
            I => \N__37269\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__37272\,
            I => \N__37266\
        );

    \I__7518\ : Odrv4
    port map (
            O => \N__37269\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__7517\ : Odrv12
    port map (
            O => \N__37266\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__7516\ : InMux
    port map (
            O => \N__37261\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__7515\ : InMux
    port map (
            O => \N__37258\,
            I => \N__37254\
        );

    \I__7514\ : CascadeMux
    port map (
            O => \N__37257\,
            I => \N__37251\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__37254\,
            I => \N__37248\
        );

    \I__7512\ : InMux
    port map (
            O => \N__37251\,
            I => \N__37245\
        );

    \I__7511\ : Span4Mux_v
    port map (
            O => \N__37248\,
            I => \N__37240\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__37245\,
            I => \N__37240\
        );

    \I__7509\ : Odrv4
    port map (
            O => \N__37240\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__7508\ : InMux
    port map (
            O => \N__37237\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__7507\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37229\
        );

    \I__7506\ : InMux
    port map (
            O => \N__37233\,
            I => \N__37226\
        );

    \I__7505\ : InMux
    port map (
            O => \N__37232\,
            I => \N__37223\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__37229\,
            I => \N__37220\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__37226\,
            I => \N__37217\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__37223\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__7501\ : Odrv4
    port map (
            O => \N__37220\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__7500\ : Odrv4
    port map (
            O => \N__37217\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__7499\ : InMux
    port map (
            O => \N__37210\,
            I => \N__37207\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__37207\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\
        );

    \I__7497\ : InMux
    port map (
            O => \N__37204\,
            I => \N__37201\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__37201\,
            I => \N__37196\
        );

    \I__7495\ : InMux
    port map (
            O => \N__37200\,
            I => \N__37193\
        );

    \I__7494\ : InMux
    port map (
            O => \N__37199\,
            I => \N__37190\
        );

    \I__7493\ : Sp12to4
    port map (
            O => \N__37196\,
            I => \N__37185\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__37193\,
            I => \N__37185\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__37190\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__7490\ : Odrv12
    port map (
            O => \N__37185\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__7489\ : InMux
    port map (
            O => \N__37180\,
            I => \N__37177\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__37177\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\
        );

    \I__7487\ : InMux
    port map (
            O => \N__37174\,
            I => \N__37169\
        );

    \I__7486\ : InMux
    port map (
            O => \N__37173\,
            I => \N__37166\
        );

    \I__7485\ : InMux
    port map (
            O => \N__37172\,
            I => \N__37163\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__37169\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__37166\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__37163\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__7481\ : CascadeMux
    port map (
            O => \N__37156\,
            I => \N__37153\
        );

    \I__7480\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37150\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__37150\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\
        );

    \I__7478\ : InMux
    port map (
            O => \N__37147\,
            I => \N__37143\
        );

    \I__7477\ : InMux
    port map (
            O => \N__37146\,
            I => \N__37140\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__37143\,
            I => \N__37137\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__37140\,
            I => \N__37134\
        );

    \I__7474\ : Span4Mux_h
    port map (
            O => \N__37137\,
            I => \N__37128\
        );

    \I__7473\ : Span4Mux_h
    port map (
            O => \N__37134\,
            I => \N__37128\
        );

    \I__7472\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37125\
        );

    \I__7471\ : Odrv4
    port map (
            O => \N__37128\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__37125\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__7469\ : CascadeMux
    port map (
            O => \N__37120\,
            I => \N__37117\
        );

    \I__7468\ : InMux
    port map (
            O => \N__37117\,
            I => \N__37112\
        );

    \I__7467\ : InMux
    port map (
            O => \N__37116\,
            I => \N__37109\
        );

    \I__7466\ : InMux
    port map (
            O => \N__37115\,
            I => \N__37106\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__37112\,
            I => \N__37103\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__37109\,
            I => \N__37100\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__37106\,
            I => \N__37095\
        );

    \I__7462\ : Span4Mux_h
    port map (
            O => \N__37103\,
            I => \N__37090\
        );

    \I__7461\ : Span4Mux_h
    port map (
            O => \N__37100\,
            I => \N__37090\
        );

    \I__7460\ : InMux
    port map (
            O => \N__37099\,
            I => \N__37085\
        );

    \I__7459\ : InMux
    port map (
            O => \N__37098\,
            I => \N__37085\
        );

    \I__7458\ : Span4Mux_h
    port map (
            O => \N__37095\,
            I => \N__37082\
        );

    \I__7457\ : Odrv4
    port map (
            O => \N__37090\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__37085\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__7455\ : Odrv4
    port map (
            O => \N__37082\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__7454\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37072\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__37072\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_20\
        );

    \I__7452\ : InMux
    port map (
            O => \N__37069\,
            I => \N__37066\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__37066\,
            I => \N__37061\
        );

    \I__7450\ : InMux
    port map (
            O => \N__37065\,
            I => \N__37058\
        );

    \I__7449\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37055\
        );

    \I__7448\ : Sp12to4
    port map (
            O => \N__37061\,
            I => \N__37050\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__37058\,
            I => \N__37050\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__37055\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__7445\ : Odrv12
    port map (
            O => \N__37050\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__7444\ : InMux
    port map (
            O => \N__37045\,
            I => \N__37042\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__37042\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\
        );

    \I__7442\ : CascadeMux
    port map (
            O => \N__37039\,
            I => \N__37036\
        );

    \I__7441\ : InMux
    port map (
            O => \N__37036\,
            I => \N__37032\
        );

    \I__7440\ : InMux
    port map (
            O => \N__37035\,
            I => \N__37028\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__37032\,
            I => \N__37025\
        );

    \I__7438\ : InMux
    port map (
            O => \N__37031\,
            I => \N__37022\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__37028\,
            I => \N__37019\
        );

    \I__7436\ : Span4Mux_v
    port map (
            O => \N__37025\,
            I => \N__37016\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__37022\,
            I => \N__37013\
        );

    \I__7434\ : Span4Mux_v
    port map (
            O => \N__37019\,
            I => \N__37010\
        );

    \I__7433\ : Span4Mux_h
    port map (
            O => \N__37016\,
            I => \N__37007\
        );

    \I__7432\ : Span4Mux_v
    port map (
            O => \N__37013\,
            I => \N__37004\
        );

    \I__7431\ : Span4Mux_h
    port map (
            O => \N__37010\,
            I => \N__37001\
        );

    \I__7430\ : Odrv4
    port map (
            O => \N__37007\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__7429\ : Odrv4
    port map (
            O => \N__37004\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__7428\ : Odrv4
    port map (
            O => \N__37001\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36994\,
            I => \N__36990\
        );

    \I__7426\ : InMux
    port map (
            O => \N__36993\,
            I => \N__36987\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__36990\,
            I => \N__36982\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__36987\,
            I => \N__36982\
        );

    \I__7423\ : Span4Mux_h
    port map (
            O => \N__36982\,
            I => \N__36979\
        );

    \I__7422\ : Odrv4
    port map (
            O => \N__36979\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__7421\ : InMux
    port map (
            O => \N__36976\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36973\,
            I => \N__36969\
        );

    \I__7419\ : InMux
    port map (
            O => \N__36972\,
            I => \N__36966\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__36969\,
            I => \N__36961\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__36966\,
            I => \N__36961\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__36961\,
            I => \N__36958\
        );

    \I__7415\ : Odrv4
    port map (
            O => \N__36958\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__7414\ : InMux
    port map (
            O => \N__36955\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__7413\ : InMux
    port map (
            O => \N__36952\,
            I => \N__36947\
        );

    \I__7412\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36942\
        );

    \I__7411\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36942\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__36947\,
            I => \N__36939\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__36942\,
            I => \N__36936\
        );

    \I__7408\ : Span4Mux_h
    port map (
            O => \N__36939\,
            I => \N__36931\
        );

    \I__7407\ : Span4Mux_h
    port map (
            O => \N__36936\,
            I => \N__36931\
        );

    \I__7406\ : Odrv4
    port map (
            O => \N__36931\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__7405\ : CascadeMux
    port map (
            O => \N__36928\,
            I => \N__36924\
        );

    \I__7404\ : CascadeMux
    port map (
            O => \N__36927\,
            I => \N__36921\
        );

    \I__7403\ : InMux
    port map (
            O => \N__36924\,
            I => \N__36918\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36921\,
            I => \N__36915\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__36918\,
            I => \N__36912\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__36915\,
            I => \N__36908\
        );

    \I__7399\ : Span4Mux_v
    port map (
            O => \N__36912\,
            I => \N__36903\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36911\,
            I => \N__36900\
        );

    \I__7397\ : Span4Mux_v
    port map (
            O => \N__36908\,
            I => \N__36897\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36907\,
            I => \N__36894\
        );

    \I__7395\ : InMux
    port map (
            O => \N__36906\,
            I => \N__36891\
        );

    \I__7394\ : Span4Mux_h
    port map (
            O => \N__36903\,
            I => \N__36886\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__36900\,
            I => \N__36886\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__36897\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__36894\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__36891\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__7389\ : Odrv4
    port map (
            O => \N__36886\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__7388\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36874\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__36874\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_19\
        );

    \I__7386\ : CascadeMux
    port map (
            O => \N__36871\,
            I => \N__36868\
        );

    \I__7385\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36865\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__36865\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_15\
        );

    \I__7383\ : InMux
    port map (
            O => \N__36862\,
            I => \N__36858\
        );

    \I__7382\ : InMux
    port map (
            O => \N__36861\,
            I => \N__36855\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__36858\,
            I => \N__36851\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__36855\,
            I => \N__36848\
        );

    \I__7379\ : InMux
    port map (
            O => \N__36854\,
            I => \N__36845\
        );

    \I__7378\ : Span4Mux_h
    port map (
            O => \N__36851\,
            I => \N__36840\
        );

    \I__7377\ : Span4Mux_h
    port map (
            O => \N__36848\,
            I => \N__36840\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__36845\,
            I => \N__36837\
        );

    \I__7375\ : Odrv4
    port map (
            O => \N__36840\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__7374\ : Odrv4
    port map (
            O => \N__36837\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__7373\ : CascadeMux
    port map (
            O => \N__36832\,
            I => \N__36828\
        );

    \I__7372\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36824\
        );

    \I__7371\ : InMux
    port map (
            O => \N__36828\,
            I => \N__36821\
        );

    \I__7370\ : InMux
    port map (
            O => \N__36827\,
            I => \N__36816\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__36824\,
            I => \N__36813\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__36821\,
            I => \N__36810\
        );

    \I__7367\ : InMux
    port map (
            O => \N__36820\,
            I => \N__36807\
        );

    \I__7366\ : CascadeMux
    port map (
            O => \N__36819\,
            I => \N__36804\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__36816\,
            I => \N__36801\
        );

    \I__7364\ : Span4Mux_v
    port map (
            O => \N__36813\,
            I => \N__36796\
        );

    \I__7363\ : Span4Mux_h
    port map (
            O => \N__36810\,
            I => \N__36796\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__36807\,
            I => \N__36793\
        );

    \I__7361\ : InMux
    port map (
            O => \N__36804\,
            I => \N__36790\
        );

    \I__7360\ : Span4Mux_h
    port map (
            O => \N__36801\,
            I => \N__36787\
        );

    \I__7359\ : Odrv4
    port map (
            O => \N__36796\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__7358\ : Odrv12
    port map (
            O => \N__36793\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__36790\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__7356\ : Odrv4
    port map (
            O => \N__36787\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__7355\ : InMux
    port map (
            O => \N__36778\,
            I => \N__36775\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__36775\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_16\
        );

    \I__7353\ : InMux
    port map (
            O => \N__36772\,
            I => \N__36768\
        );

    \I__7352\ : InMux
    port map (
            O => \N__36771\,
            I => \N__36765\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__36768\,
            I => \N__36761\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__36765\,
            I => \N__36758\
        );

    \I__7349\ : InMux
    port map (
            O => \N__36764\,
            I => \N__36755\
        );

    \I__7348\ : Span4Mux_h
    port map (
            O => \N__36761\,
            I => \N__36752\
        );

    \I__7347\ : Span4Mux_h
    port map (
            O => \N__36758\,
            I => \N__36749\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__36755\,
            I => \N__36746\
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__36752\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__36749\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__7343\ : Odrv4
    port map (
            O => \N__36746\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__7342\ : InMux
    port map (
            O => \N__36739\,
            I => \N__36735\
        );

    \I__7341\ : InMux
    port map (
            O => \N__36738\,
            I => \N__36732\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__36735\,
            I => \N__36729\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__36732\,
            I => \N__36726\
        );

    \I__7338\ : Span4Mux_h
    port map (
            O => \N__36729\,
            I => \N__36722\
        );

    \I__7337\ : Span4Mux_h
    port map (
            O => \N__36726\,
            I => \N__36719\
        );

    \I__7336\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36716\
        );

    \I__7335\ : Odrv4
    port map (
            O => \N__36722\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__7334\ : Odrv4
    port map (
            O => \N__36719\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__36716\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__7332\ : InMux
    port map (
            O => \N__36709\,
            I => \N__36706\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__36706\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_23\
        );

    \I__7330\ : InMux
    port map (
            O => \N__36703\,
            I => \N__36699\
        );

    \I__7329\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36696\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__36699\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__36696\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__7326\ : CascadeMux
    port map (
            O => \N__36691\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_\
        );

    \I__7325\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36685\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__36685\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\
        );

    \I__7323\ : InMux
    port map (
            O => \N__36682\,
            I => \N__36679\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__36679\,
            I => \N__36674\
        );

    \I__7321\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36671\
        );

    \I__7320\ : InMux
    port map (
            O => \N__36677\,
            I => \N__36668\
        );

    \I__7319\ : Span4Mux_h
    port map (
            O => \N__36674\,
            I => \N__36665\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__36671\,
            I => \N__36660\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__36668\,
            I => \N__36660\
        );

    \I__7316\ : Odrv4
    port map (
            O => \N__36665\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__7315\ : Odrv4
    port map (
            O => \N__36660\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__7314\ : InMux
    port map (
            O => \N__36655\,
            I => \N__36652\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__36652\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_7\
        );

    \I__7312\ : CascadeMux
    port map (
            O => \N__36649\,
            I => \N__36646\
        );

    \I__7311\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36643\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__36643\,
            I => \N__36639\
        );

    \I__7309\ : InMux
    port map (
            O => \N__36642\,
            I => \N__36635\
        );

    \I__7308\ : Span4Mux_h
    port map (
            O => \N__36639\,
            I => \N__36632\
        );

    \I__7307\ : InMux
    port map (
            O => \N__36638\,
            I => \N__36629\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__36635\,
            I => \N__36626\
        );

    \I__7305\ : Span4Mux_h
    port map (
            O => \N__36632\,
            I => \N__36621\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__36629\,
            I => \N__36621\
        );

    \I__7303\ : Odrv12
    port map (
            O => \N__36626\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__7302\ : Odrv4
    port map (
            O => \N__36621\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__7301\ : InMux
    port map (
            O => \N__36616\,
            I => \N__36613\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__36613\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_9\
        );

    \I__7299\ : InMux
    port map (
            O => \N__36610\,
            I => \N__36606\
        );

    \I__7298\ : InMux
    port map (
            O => \N__36609\,
            I => \N__36603\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__36606\,
            I => \N__36599\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__36603\,
            I => \N__36596\
        );

    \I__7295\ : InMux
    port map (
            O => \N__36602\,
            I => \N__36593\
        );

    \I__7294\ : Span4Mux_h
    port map (
            O => \N__36599\,
            I => \N__36590\
        );

    \I__7293\ : Span4Mux_h
    port map (
            O => \N__36596\,
            I => \N__36585\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__36593\,
            I => \N__36585\
        );

    \I__7291\ : Odrv4
    port map (
            O => \N__36590\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__7290\ : Odrv4
    port map (
            O => \N__36585\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__7289\ : InMux
    port map (
            O => \N__36580\,
            I => \N__36577\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__36577\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_10\
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__36574\,
            I => \N__36571\
        );

    \I__7286\ : InMux
    port map (
            O => \N__36571\,
            I => \N__36567\
        );

    \I__7285\ : InMux
    port map (
            O => \N__36570\,
            I => \N__36564\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__36567\,
            I => \N__36561\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__36564\,
            I => \N__36557\
        );

    \I__7282\ : Span4Mux_v
    port map (
            O => \N__36561\,
            I => \N__36554\
        );

    \I__7281\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36551\
        );

    \I__7280\ : Span4Mux_v
    port map (
            O => \N__36557\,
            I => \N__36546\
        );

    \I__7279\ : Span4Mux_v
    port map (
            O => \N__36554\,
            I => \N__36546\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__36551\,
            I => \N__36543\
        );

    \I__7277\ : Odrv4
    port map (
            O => \N__36546\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7276\ : Odrv4
    port map (
            O => \N__36543\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7275\ : InMux
    port map (
            O => \N__36538\,
            I => \N__36535\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__36535\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_12\
        );

    \I__7273\ : CascadeMux
    port map (
            O => \N__36532\,
            I => \N__36527\
        );

    \I__7272\ : InMux
    port map (
            O => \N__36531\,
            I => \N__36524\
        );

    \I__7271\ : InMux
    port map (
            O => \N__36530\,
            I => \N__36521\
        );

    \I__7270\ : InMux
    port map (
            O => \N__36527\,
            I => \N__36518\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__36524\,
            I => \N__36514\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__36521\,
            I => \N__36511\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__36518\,
            I => \N__36508\
        );

    \I__7266\ : InMux
    port map (
            O => \N__36517\,
            I => \N__36505\
        );

    \I__7265\ : Span4Mux_v
    port map (
            O => \N__36514\,
            I => \N__36502\
        );

    \I__7264\ : Span4Mux_v
    port map (
            O => \N__36511\,
            I => \N__36499\
        );

    \I__7263\ : Span4Mux_h
    port map (
            O => \N__36508\,
            I => \N__36492\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__36505\,
            I => \N__36492\
        );

    \I__7261\ : Span4Mux_h
    port map (
            O => \N__36502\,
            I => \N__36492\
        );

    \I__7260\ : Odrv4
    port map (
            O => \N__36499\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__7259\ : Odrv4
    port map (
            O => \N__36492\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__7258\ : InMux
    port map (
            O => \N__36487\,
            I => \N__36483\
        );

    \I__7257\ : InMux
    port map (
            O => \N__36486\,
            I => \N__36480\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__36483\,
            I => \N__36476\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__36480\,
            I => \N__36473\
        );

    \I__7254\ : InMux
    port map (
            O => \N__36479\,
            I => \N__36470\
        );

    \I__7253\ : Span4Mux_h
    port map (
            O => \N__36476\,
            I => \N__36465\
        );

    \I__7252\ : Span4Mux_v
    port map (
            O => \N__36473\,
            I => \N__36465\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__36470\,
            I => \N__36462\
        );

    \I__7250\ : Odrv4
    port map (
            O => \N__36465\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__7249\ : Odrv4
    port map (
            O => \N__36462\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__7248\ : InMux
    port map (
            O => \N__36457\,
            I => \N__36454\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__36454\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_11\
        );

    \I__7246\ : InMux
    port map (
            O => \N__36451\,
            I => \N__36447\
        );

    \I__7245\ : InMux
    port map (
            O => \N__36450\,
            I => \N__36444\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__36447\,
            I => \N__36441\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__36444\,
            I => \N__36438\
        );

    \I__7242\ : Span4Mux_h
    port map (
            O => \N__36441\,
            I => \N__36434\
        );

    \I__7241\ : Span4Mux_h
    port map (
            O => \N__36438\,
            I => \N__36431\
        );

    \I__7240\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36428\
        );

    \I__7239\ : Odrv4
    port map (
            O => \N__36434\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__36431\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__36428\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__7236\ : InMux
    port map (
            O => \N__36421\,
            I => \N__36418\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__36418\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_22\
        );

    \I__7234\ : CEMux
    port map (
            O => \N__36415\,
            I => \N__36412\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__36412\,
            I => \N__36406\
        );

    \I__7232\ : CEMux
    port map (
            O => \N__36411\,
            I => \N__36403\
        );

    \I__7231\ : CEMux
    port map (
            O => \N__36410\,
            I => \N__36400\
        );

    \I__7230\ : CEMux
    port map (
            O => \N__36409\,
            I => \N__36396\
        );

    \I__7229\ : Span4Mux_h
    port map (
            O => \N__36406\,
            I => \N__36392\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__36403\,
            I => \N__36389\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__36400\,
            I => \N__36386\
        );

    \I__7226\ : CEMux
    port map (
            O => \N__36399\,
            I => \N__36383\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__36396\,
            I => \N__36380\
        );

    \I__7224\ : IoInMux
    port map (
            O => \N__36395\,
            I => \N__36377\
        );

    \I__7223\ : Sp12to4
    port map (
            O => \N__36392\,
            I => \N__36374\
        );

    \I__7222\ : Span4Mux_v
    port map (
            O => \N__36389\,
            I => \N__36371\
        );

    \I__7221\ : Span4Mux_h
    port map (
            O => \N__36386\,
            I => \N__36366\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__36383\,
            I => \N__36366\
        );

    \I__7219\ : Span4Mux_v
    port map (
            O => \N__36380\,
            I => \N__36363\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__36377\,
            I => \N__36360\
        );

    \I__7217\ : Span12Mux_v
    port map (
            O => \N__36374\,
            I => \N__36357\
        );

    \I__7216\ : Sp12to4
    port map (
            O => \N__36371\,
            I => \N__36354\
        );

    \I__7215\ : Span4Mux_v
    port map (
            O => \N__36366\,
            I => \N__36351\
        );

    \I__7214\ : Span4Mux_v
    port map (
            O => \N__36363\,
            I => \N__36348\
        );

    \I__7213\ : Span4Mux_s2_v
    port map (
            O => \N__36360\,
            I => \N__36345\
        );

    \I__7212\ : Span12Mux_v
    port map (
            O => \N__36357\,
            I => \N__36342\
        );

    \I__7211\ : Span12Mux_v
    port map (
            O => \N__36354\,
            I => \N__36339\
        );

    \I__7210\ : Span4Mux_v
    port map (
            O => \N__36351\,
            I => \N__36336\
        );

    \I__7209\ : Span4Mux_v
    port map (
            O => \N__36348\,
            I => \N__36331\
        );

    \I__7208\ : Span4Mux_h
    port map (
            O => \N__36345\,
            I => \N__36331\
        );

    \I__7207\ : Odrv12
    port map (
            O => \N__36342\,
            I => red_c_i
        );

    \I__7206\ : Odrv12
    port map (
            O => \N__36339\,
            I => red_c_i
        );

    \I__7205\ : Odrv4
    port map (
            O => \N__36336\,
            I => red_c_i
        );

    \I__7204\ : Odrv4
    port map (
            O => \N__36331\,
            I => red_c_i
        );

    \I__7203\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36318\
        );

    \I__7202\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36315\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__36318\,
            I => \N__36312\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__36315\,
            I => \N__36308\
        );

    \I__7199\ : Span4Mux_h
    port map (
            O => \N__36312\,
            I => \N__36305\
        );

    \I__7198\ : InMux
    port map (
            O => \N__36311\,
            I => \N__36302\
        );

    \I__7197\ : Span4Mux_h
    port map (
            O => \N__36308\,
            I => \N__36299\
        );

    \I__7196\ : Span4Mux_v
    port map (
            O => \N__36305\,
            I => \N__36296\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__36302\,
            I => \N__36293\
        );

    \I__7194\ : Odrv4
    port map (
            O => \N__36299\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__7193\ : Odrv4
    port map (
            O => \N__36296\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__7192\ : Odrv4
    port map (
            O => \N__36293\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__7191\ : InMux
    port map (
            O => \N__36286\,
            I => \N__36283\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__36283\,
            I => \N__36280\
        );

    \I__7189\ : Odrv4
    port map (
            O => \N__36280\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_13\
        );

    \I__7188\ : InMux
    port map (
            O => \N__36277\,
            I => \N__36273\
        );

    \I__7187\ : InMux
    port map (
            O => \N__36276\,
            I => \N__36270\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__36273\,
            I => \N__36266\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__36270\,
            I => \N__36263\
        );

    \I__7184\ : InMux
    port map (
            O => \N__36269\,
            I => \N__36260\
        );

    \I__7183\ : Span4Mux_h
    port map (
            O => \N__36266\,
            I => \N__36257\
        );

    \I__7182\ : Span4Mux_h
    port map (
            O => \N__36263\,
            I => \N__36252\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__36260\,
            I => \N__36252\
        );

    \I__7180\ : Odrv4
    port map (
            O => \N__36257\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__7179\ : Odrv4
    port map (
            O => \N__36252\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__7178\ : InMux
    port map (
            O => \N__36247\,
            I => \N__36244\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__36244\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_6\
        );

    \I__7176\ : InMux
    port map (
            O => \N__36241\,
            I => \N__36237\
        );

    \I__7175\ : InMux
    port map (
            O => \N__36240\,
            I => \N__36234\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__36237\,
            I => \N__36230\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__36234\,
            I => \N__36227\
        );

    \I__7172\ : InMux
    port map (
            O => \N__36233\,
            I => \N__36224\
        );

    \I__7171\ : Span4Mux_v
    port map (
            O => \N__36230\,
            I => \N__36219\
        );

    \I__7170\ : Span4Mux_v
    port map (
            O => \N__36227\,
            I => \N__36219\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__36224\,
            I => \N__36216\
        );

    \I__7168\ : Odrv4
    port map (
            O => \N__36219\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__7167\ : Odrv4
    port map (
            O => \N__36216\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__7166\ : InMux
    port map (
            O => \N__36211\,
            I => \N__36208\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__36208\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_5\
        );

    \I__7164\ : InMux
    port map (
            O => \N__36205\,
            I => \N__36201\
        );

    \I__7163\ : InMux
    port map (
            O => \N__36204\,
            I => \N__36198\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__36201\,
            I => \N__36194\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__36198\,
            I => \N__36191\
        );

    \I__7160\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36188\
        );

    \I__7159\ : Span4Mux_v
    port map (
            O => \N__36194\,
            I => \N__36183\
        );

    \I__7158\ : Span4Mux_v
    port map (
            O => \N__36191\,
            I => \N__36183\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__36188\,
            I => \N__36180\
        );

    \I__7156\ : Odrv4
    port map (
            O => \N__36183\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__7155\ : Odrv4
    port map (
            O => \N__36180\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__7154\ : InMux
    port map (
            O => \N__36175\,
            I => \N__36172\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__36172\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_4\
        );

    \I__7152\ : InMux
    port map (
            O => \N__36169\,
            I => \N__36165\
        );

    \I__7151\ : InMux
    port map (
            O => \N__36168\,
            I => \N__36162\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__36165\,
            I => \N__36158\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__36162\,
            I => \N__36155\
        );

    \I__7148\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36152\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__36158\,
            I => \N__36149\
        );

    \I__7146\ : Span4Mux_h
    port map (
            O => \N__36155\,
            I => \N__36144\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__36152\,
            I => \N__36144\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__36149\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__36144\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__7142\ : InMux
    port map (
            O => \N__36139\,
            I => \N__36136\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__36136\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_8\
        );

    \I__7140\ : InMux
    port map (
            O => \N__36133\,
            I => \N__36127\
        );

    \I__7139\ : InMux
    port map (
            O => \N__36132\,
            I => \N__36127\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__36127\,
            I => \N__36123\
        );

    \I__7137\ : InMux
    port map (
            O => \N__36126\,
            I => \N__36120\
        );

    \I__7136\ : Span4Mux_v
    port map (
            O => \N__36123\,
            I => \N__36117\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__36120\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__36117\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__7133\ : CascadeMux
    port map (
            O => \N__36112\,
            I => \N__36109\
        );

    \I__7132\ : InMux
    port map (
            O => \N__36109\,
            I => \N__36106\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__36106\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__7130\ : InMux
    port map (
            O => \N__36103\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__7129\ : CascadeMux
    port map (
            O => \N__36100\,
            I => \N__36096\
        );

    \I__7128\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36093\
        );

    \I__7127\ : InMux
    port map (
            O => \N__36096\,
            I => \N__36090\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__36093\,
            I => \N__36084\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__36090\,
            I => \N__36084\
        );

    \I__7124\ : InMux
    port map (
            O => \N__36089\,
            I => \N__36081\
        );

    \I__7123\ : Span4Mux_v
    port map (
            O => \N__36084\,
            I => \N__36078\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__36081\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__36078\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__7120\ : InMux
    port map (
            O => \N__36073\,
            I => \N__36070\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__36070\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__7118\ : InMux
    port map (
            O => \N__36067\,
            I => \bfn_14_29_0_\
        );

    \I__7117\ : InMux
    port map (
            O => \N__36064\,
            I => \N__36060\
        );

    \I__7116\ : CascadeMux
    port map (
            O => \N__36063\,
            I => \N__36057\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__36060\,
            I => \N__36054\
        );

    \I__7114\ : InMux
    port map (
            O => \N__36057\,
            I => \N__36051\
        );

    \I__7113\ : Span4Mux_s2_v
    port map (
            O => \N__36054\,
            I => \N__36045\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__36051\,
            I => \N__36045\
        );

    \I__7111\ : InMux
    port map (
            O => \N__36050\,
            I => \N__36042\
        );

    \I__7110\ : Span4Mux_v
    port map (
            O => \N__36045\,
            I => \N__36039\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__36042\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__7108\ : Odrv4
    port map (
            O => \N__36039\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__7107\ : InMux
    port map (
            O => \N__36034\,
            I => \N__36031\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__36031\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__7105\ : InMux
    port map (
            O => \N__36028\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__7104\ : CascadeMux
    port map (
            O => \N__36025\,
            I => \N__36021\
        );

    \I__7103\ : InMux
    port map (
            O => \N__36024\,
            I => \N__36017\
        );

    \I__7102\ : InMux
    port map (
            O => \N__36021\,
            I => \N__36014\
        );

    \I__7101\ : InMux
    port map (
            O => \N__36020\,
            I => \N__36011\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__36017\,
            I => \N__36006\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__36014\,
            I => \N__36006\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__36011\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__7097\ : Odrv12
    port map (
            O => \N__36006\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__36001\,
            I => \N__35998\
        );

    \I__7095\ : InMux
    port map (
            O => \N__35998\,
            I => \N__35995\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__35995\,
            I => \N__35991\
        );

    \I__7093\ : InMux
    port map (
            O => \N__35994\,
            I => \N__35988\
        );

    \I__7092\ : Span4Mux_s3_v
    port map (
            O => \N__35991\,
            I => \N__35985\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__35988\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__7090\ : Odrv4
    port map (
            O => \N__35985\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__7089\ : InMux
    port map (
            O => \N__35980\,
            I => \N__35977\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__35977\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35974\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__7086\ : CascadeMux
    port map (
            O => \N__35971\,
            I => \N__35967\
        );

    \I__7085\ : InMux
    port map (
            O => \N__35970\,
            I => \N__35963\
        );

    \I__7084\ : InMux
    port map (
            O => \N__35967\,
            I => \N__35960\
        );

    \I__7083\ : InMux
    port map (
            O => \N__35966\,
            I => \N__35957\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__35963\,
            I => \N__35952\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__35960\,
            I => \N__35952\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__35957\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__7079\ : Odrv12
    port map (
            O => \N__35952\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__7078\ : CascadeMux
    port map (
            O => \N__35947\,
            I => \N__35944\
        );

    \I__7077\ : InMux
    port map (
            O => \N__35944\,
            I => \N__35940\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35943\,
            I => \N__35937\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__35940\,
            I => \N__35934\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__35937\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__7073\ : Odrv12
    port map (
            O => \N__35934\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__7072\ : CascadeMux
    port map (
            O => \N__35929\,
            I => \N__35926\
        );

    \I__7071\ : InMux
    port map (
            O => \N__35926\,
            I => \N__35923\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__35923\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__7069\ : InMux
    port map (
            O => \N__35920\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__7068\ : InMux
    port map (
            O => \N__35917\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__7067\ : InMux
    port map (
            O => \N__35914\,
            I => \N__35911\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__35911\,
            I => \N__35907\
        );

    \I__7065\ : InMux
    port map (
            O => \N__35910\,
            I => \N__35904\
        );

    \I__7064\ : Odrv4
    port map (
            O => \N__35907\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__35904\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__7062\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35896\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__35896\,
            I => \N__35893\
        );

    \I__7060\ : Odrv12
    port map (
            O => \N__35893\,
            I => delay_tr_input_c
        );

    \I__7059\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35887\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__35887\,
            I => delay_tr_d1
        );

    \I__7057\ : InMux
    port map (
            O => \N__35884\,
            I => \N__35878\
        );

    \I__7056\ : InMux
    port map (
            O => \N__35883\,
            I => \N__35878\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__35878\,
            I => \N__35874\
        );

    \I__7054\ : InMux
    port map (
            O => \N__35877\,
            I => \N__35871\
        );

    \I__7053\ : Span4Mux_v
    port map (
            O => \N__35874\,
            I => \N__35868\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__35871\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__7051\ : Odrv4
    port map (
            O => \N__35868\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__7050\ : InMux
    port map (
            O => \N__35863\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__7049\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35856\
        );

    \I__7048\ : CascadeMux
    port map (
            O => \N__35859\,
            I => \N__35853\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__35856\,
            I => \N__35850\
        );

    \I__7046\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35847\
        );

    \I__7045\ : Span4Mux_s3_v
    port map (
            O => \N__35850\,
            I => \N__35841\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__35847\,
            I => \N__35841\
        );

    \I__7043\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35838\
        );

    \I__7042\ : Span4Mux_v
    port map (
            O => \N__35841\,
            I => \N__35835\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__35838\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__7040\ : Odrv4
    port map (
            O => \N__35835\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__7039\ : InMux
    port map (
            O => \N__35830\,
            I => \bfn_14_28_0_\
        );

    \I__7038\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35823\
        );

    \I__7037\ : CascadeMux
    port map (
            O => \N__35826\,
            I => \N__35820\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__35823\,
            I => \N__35817\
        );

    \I__7035\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35814\
        );

    \I__7034\ : Span4Mux_s3_v
    port map (
            O => \N__35817\,
            I => \N__35808\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__35814\,
            I => \N__35808\
        );

    \I__7032\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35805\
        );

    \I__7031\ : Span4Mux_v
    port map (
            O => \N__35808\,
            I => \N__35802\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__35805\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__35802\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__7028\ : CascadeMux
    port map (
            O => \N__35797\,
            I => \N__35793\
        );

    \I__7027\ : InMux
    port map (
            O => \N__35796\,
            I => \N__35790\
        );

    \I__7026\ : InMux
    port map (
            O => \N__35793\,
            I => \N__35787\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__35790\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__35787\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__7023\ : InMux
    port map (
            O => \N__35782\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__7022\ : CascadeMux
    port map (
            O => \N__35779\,
            I => \N__35775\
        );

    \I__7021\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35771\
        );

    \I__7020\ : InMux
    port map (
            O => \N__35775\,
            I => \N__35768\
        );

    \I__7019\ : InMux
    port map (
            O => \N__35774\,
            I => \N__35765\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__35771\,
            I => \N__35760\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__35768\,
            I => \N__35760\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__35765\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__7015\ : Odrv12
    port map (
            O => \N__35760\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__7014\ : InMux
    port map (
            O => \N__35755\,
            I => \N__35749\
        );

    \I__7013\ : InMux
    port map (
            O => \N__35754\,
            I => \N__35749\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__35749\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__7011\ : InMux
    port map (
            O => \N__35746\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__7010\ : CascadeMux
    port map (
            O => \N__35743\,
            I => \N__35739\
        );

    \I__7009\ : InMux
    port map (
            O => \N__35742\,
            I => \N__35735\
        );

    \I__7008\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35732\
        );

    \I__7007\ : InMux
    port map (
            O => \N__35738\,
            I => \N__35729\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__35735\,
            I => \N__35724\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__35732\,
            I => \N__35724\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__35729\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__7003\ : Odrv12
    port map (
            O => \N__35724\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__7002\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35713\
        );

    \I__7001\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35713\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__35713\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__6999\ : InMux
    port map (
            O => \N__35710\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__6998\ : CascadeMux
    port map (
            O => \N__35707\,
            I => \N__35703\
        );

    \I__6997\ : CascadeMux
    port map (
            O => \N__35706\,
            I => \N__35700\
        );

    \I__6996\ : InMux
    port map (
            O => \N__35703\,
            I => \N__35695\
        );

    \I__6995\ : InMux
    port map (
            O => \N__35700\,
            I => \N__35695\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__35695\,
            I => \N__35691\
        );

    \I__6993\ : InMux
    port map (
            O => \N__35694\,
            I => \N__35688\
        );

    \I__6992\ : Span4Mux_v
    port map (
            O => \N__35691\,
            I => \N__35685\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__35688\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__6990\ : Odrv4
    port map (
            O => \N__35685\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__6989\ : InMux
    port map (
            O => \N__35680\,
            I => \N__35677\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__35677\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__6987\ : InMux
    port map (
            O => \N__35674\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__6986\ : CascadeMux
    port map (
            O => \N__35671\,
            I => \N__35667\
        );

    \I__6985\ : CascadeMux
    port map (
            O => \N__35670\,
            I => \N__35664\
        );

    \I__6984\ : InMux
    port map (
            O => \N__35667\,
            I => \N__35658\
        );

    \I__6983\ : InMux
    port map (
            O => \N__35664\,
            I => \N__35658\
        );

    \I__6982\ : InMux
    port map (
            O => \N__35663\,
            I => \N__35655\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__35658\,
            I => \N__35652\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__35655\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__6979\ : Odrv12
    port map (
            O => \N__35652\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__6978\ : InMux
    port map (
            O => \N__35647\,
            I => \N__35644\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__35644\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__6976\ : InMux
    port map (
            O => \N__35641\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__6975\ : InMux
    port map (
            O => \N__35638\,
            I => \N__35632\
        );

    \I__6974\ : InMux
    port map (
            O => \N__35637\,
            I => \N__35632\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__35632\,
            I => \N__35628\
        );

    \I__6972\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35625\
        );

    \I__6971\ : Span4Mux_v
    port map (
            O => \N__35628\,
            I => \N__35622\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__35625\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__6969\ : Odrv4
    port map (
            O => \N__35622\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__6968\ : InMux
    port map (
            O => \N__35617\,
            I => \N__35614\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__35614\,
            I => \N__35611\
        );

    \I__6966\ : Odrv4
    port map (
            O => \N__35611\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__6965\ : InMux
    port map (
            O => \N__35608\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__6964\ : CascadeMux
    port map (
            O => \N__35605\,
            I => \N__35601\
        );

    \I__6963\ : CascadeMux
    port map (
            O => \N__35604\,
            I => \N__35598\
        );

    \I__6962\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35593\
        );

    \I__6961\ : InMux
    port map (
            O => \N__35598\,
            I => \N__35593\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__35593\,
            I => \N__35589\
        );

    \I__6959\ : InMux
    port map (
            O => \N__35592\,
            I => \N__35586\
        );

    \I__6958\ : Span4Mux_v
    port map (
            O => \N__35589\,
            I => \N__35583\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__35586\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__6956\ : Odrv4
    port map (
            O => \N__35583\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__6955\ : InMux
    port map (
            O => \N__35578\,
            I => \N__35574\
        );

    \I__6954\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35571\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__35574\,
            I => \N__35568\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__35571\,
            I => \N__35565\
        );

    \I__6951\ : Span4Mux_h
    port map (
            O => \N__35568\,
            I => \N__35561\
        );

    \I__6950\ : Span4Mux_h
    port map (
            O => \N__35565\,
            I => \N__35558\
        );

    \I__6949\ : InMux
    port map (
            O => \N__35564\,
            I => \N__35555\
        );

    \I__6948\ : Odrv4
    port map (
            O => \N__35561\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__6947\ : Odrv4
    port map (
            O => \N__35558\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__35555\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__6945\ : InMux
    port map (
            O => \N__35548\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__6944\ : CascadeMux
    port map (
            O => \N__35545\,
            I => \N__35541\
        );

    \I__6943\ : InMux
    port map (
            O => \N__35544\,
            I => \N__35537\
        );

    \I__6942\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35534\
        );

    \I__6941\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35531\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__35537\,
            I => \N__35526\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__35534\,
            I => \N__35526\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__35531\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__6937\ : Odrv12
    port map (
            O => \N__35526\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__6936\ : InMux
    port map (
            O => \N__35521\,
            I => \N__35518\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__35518\,
            I => \N__35513\
        );

    \I__6934\ : InMux
    port map (
            O => \N__35517\,
            I => \N__35510\
        );

    \I__6933\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35507\
        );

    \I__6932\ : Span4Mux_v
    port map (
            O => \N__35513\,
            I => \N__35502\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__35510\,
            I => \N__35502\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__35507\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__35502\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__6928\ : InMux
    port map (
            O => \N__35497\,
            I => \bfn_14_27_0_\
        );

    \I__6927\ : InMux
    port map (
            O => \N__35494\,
            I => \N__35491\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__35491\,
            I => \N__35487\
        );

    \I__6925\ : InMux
    port map (
            O => \N__35490\,
            I => \N__35484\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__35487\,
            I => \N__35478\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__35484\,
            I => \N__35478\
        );

    \I__6922\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35475\
        );

    \I__6921\ : Span4Mux_v
    port map (
            O => \N__35478\,
            I => \N__35472\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__35475\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__6919\ : Odrv4
    port map (
            O => \N__35472\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__6918\ : InMux
    port map (
            O => \N__35467\,
            I => \N__35463\
        );

    \I__6917\ : InMux
    port map (
            O => \N__35466\,
            I => \N__35460\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__35463\,
            I => \N__35456\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__35460\,
            I => \N__35453\
        );

    \I__6914\ : InMux
    port map (
            O => \N__35459\,
            I => \N__35450\
        );

    \I__6913\ : Span4Mux_v
    port map (
            O => \N__35456\,
            I => \N__35445\
        );

    \I__6912\ : Span4Mux_h
    port map (
            O => \N__35453\,
            I => \N__35445\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__35450\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__6910\ : Odrv4
    port map (
            O => \N__35445\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__6909\ : InMux
    port map (
            O => \N__35440\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__6908\ : CascadeMux
    port map (
            O => \N__35437\,
            I => \N__35433\
        );

    \I__6907\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35429\
        );

    \I__6906\ : InMux
    port map (
            O => \N__35433\,
            I => \N__35426\
        );

    \I__6905\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35423\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__35429\,
            I => \N__35418\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__35426\,
            I => \N__35418\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__35423\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__6901\ : Odrv12
    port map (
            O => \N__35418\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__6900\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35409\
        );

    \I__6899\ : CascadeMux
    port map (
            O => \N__35412\,
            I => \N__35406\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__35409\,
            I => \N__35403\
        );

    \I__6897\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35399\
        );

    \I__6896\ : Span4Mux_h
    port map (
            O => \N__35403\,
            I => \N__35396\
        );

    \I__6895\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35393\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__35399\,
            I => \N__35390\
        );

    \I__6893\ : Odrv4
    port map (
            O => \N__35396\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__35393\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__6891\ : Odrv4
    port map (
            O => \N__35390\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__6890\ : InMux
    port map (
            O => \N__35383\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__6889\ : CascadeMux
    port map (
            O => \N__35380\,
            I => \N__35376\
        );

    \I__6888\ : InMux
    port map (
            O => \N__35379\,
            I => \N__35372\
        );

    \I__6887\ : InMux
    port map (
            O => \N__35376\,
            I => \N__35369\
        );

    \I__6886\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35366\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__35372\,
            I => \N__35361\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__35369\,
            I => \N__35361\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__35366\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__6882\ : Odrv12
    port map (
            O => \N__35361\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__6881\ : InMux
    port map (
            O => \N__35356\,
            I => \N__35353\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__35353\,
            I => \N__35350\
        );

    \I__6879\ : Span4Mux_h
    port map (
            O => \N__35350\,
            I => \N__35344\
        );

    \I__6878\ : InMux
    port map (
            O => \N__35349\,
            I => \N__35339\
        );

    \I__6877\ : InMux
    port map (
            O => \N__35348\,
            I => \N__35339\
        );

    \I__6876\ : InMux
    port map (
            O => \N__35347\,
            I => \N__35336\
        );

    \I__6875\ : Odrv4
    port map (
            O => \N__35344\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__35339\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__35336\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__6872\ : InMux
    port map (
            O => \N__35329\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__6871\ : CascadeMux
    port map (
            O => \N__35326\,
            I => \N__35322\
        );

    \I__6870\ : CascadeMux
    port map (
            O => \N__35325\,
            I => \N__35319\
        );

    \I__6869\ : InMux
    port map (
            O => \N__35322\,
            I => \N__35314\
        );

    \I__6868\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35314\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__35314\,
            I => \N__35310\
        );

    \I__6866\ : InMux
    port map (
            O => \N__35313\,
            I => \N__35307\
        );

    \I__6865\ : Span4Mux_v
    port map (
            O => \N__35310\,
            I => \N__35304\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__35307\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__35304\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__6862\ : InMux
    port map (
            O => \N__35299\,
            I => \N__35295\
        );

    \I__6861\ : CascadeMux
    port map (
            O => \N__35298\,
            I => \N__35290\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__35295\,
            I => \N__35287\
        );

    \I__6859\ : InMux
    port map (
            O => \N__35294\,
            I => \N__35284\
        );

    \I__6858\ : InMux
    port map (
            O => \N__35293\,
            I => \N__35279\
        );

    \I__6857\ : InMux
    port map (
            O => \N__35290\,
            I => \N__35279\
        );

    \I__6856\ : Odrv4
    port map (
            O => \N__35287\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__35284\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__35279\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__6853\ : InMux
    port map (
            O => \N__35272\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__6852\ : CascadeMux
    port map (
            O => \N__35269\,
            I => \N__35265\
        );

    \I__6851\ : CascadeMux
    port map (
            O => \N__35268\,
            I => \N__35262\
        );

    \I__6850\ : InMux
    port map (
            O => \N__35265\,
            I => \N__35256\
        );

    \I__6849\ : InMux
    port map (
            O => \N__35262\,
            I => \N__35256\
        );

    \I__6848\ : InMux
    port map (
            O => \N__35261\,
            I => \N__35253\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__35256\,
            I => \N__35250\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__35253\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__6845\ : Odrv12
    port map (
            O => \N__35250\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__6844\ : InMux
    port map (
            O => \N__35245\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__6843\ : InMux
    port map (
            O => \N__35242\,
            I => \N__35236\
        );

    \I__6842\ : InMux
    port map (
            O => \N__35241\,
            I => \N__35236\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__35236\,
            I => \N__35232\
        );

    \I__6840\ : InMux
    port map (
            O => \N__35235\,
            I => \N__35229\
        );

    \I__6839\ : Span4Mux_v
    port map (
            O => \N__35232\,
            I => \N__35226\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__35229\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__35226\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__6836\ : InMux
    port map (
            O => \N__35221\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__6835\ : CascadeMux
    port map (
            O => \N__35218\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_\
        );

    \I__6834\ : InMux
    port map (
            O => \N__35215\,
            I => \N__35212\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__35212\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_10\
        );

    \I__6832\ : InMux
    port map (
            O => \N__35209\,
            I => \N__35206\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__35206\,
            I => \N__35203\
        );

    \I__6830\ : Span4Mux_h
    port map (
            O => \N__35203\,
            I => \N__35198\
        );

    \I__6829\ : InMux
    port map (
            O => \N__35202\,
            I => \N__35195\
        );

    \I__6828\ : InMux
    port map (
            O => \N__35201\,
            I => \N__35192\
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__35198\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__35195\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__35192\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__6824\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35180\
        );

    \I__6823\ : InMux
    port map (
            O => \N__35184\,
            I => \N__35175\
        );

    \I__6822\ : InMux
    port map (
            O => \N__35183\,
            I => \N__35175\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__35180\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__35175\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__6819\ : InMux
    port map (
            O => \N__35170\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__6818\ : CascadeMux
    port map (
            O => \N__35167\,
            I => \N__35163\
        );

    \I__6817\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35159\
        );

    \I__6816\ : InMux
    port map (
            O => \N__35163\,
            I => \N__35156\
        );

    \I__6815\ : InMux
    port map (
            O => \N__35162\,
            I => \N__35153\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__35159\,
            I => \N__35148\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__35156\,
            I => \N__35148\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__35153\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__6811\ : Odrv12
    port map (
            O => \N__35148\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__6810\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35140\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__35140\,
            I => \N__35137\
        );

    \I__6808\ : Span4Mux_h
    port map (
            O => \N__35137\,
            I => \N__35132\
        );

    \I__6807\ : InMux
    port map (
            O => \N__35136\,
            I => \N__35127\
        );

    \I__6806\ : InMux
    port map (
            O => \N__35135\,
            I => \N__35127\
        );

    \I__6805\ : Odrv4
    port map (
            O => \N__35132\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__35127\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__6803\ : InMux
    port map (
            O => \N__35122\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__6802\ : CascadeMux
    port map (
            O => \N__35119\,
            I => \N__35115\
        );

    \I__6801\ : InMux
    port map (
            O => \N__35118\,
            I => \N__35111\
        );

    \I__6800\ : InMux
    port map (
            O => \N__35115\,
            I => \N__35108\
        );

    \I__6799\ : InMux
    port map (
            O => \N__35114\,
            I => \N__35105\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__35111\,
            I => \N__35100\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__35108\,
            I => \N__35100\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__35105\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__6795\ : Odrv12
    port map (
            O => \N__35100\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__6794\ : InMux
    port map (
            O => \N__35095\,
            I => \N__35092\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__35092\,
            I => \N__35086\
        );

    \I__6792\ : InMux
    port map (
            O => \N__35091\,
            I => \N__35079\
        );

    \I__6791\ : InMux
    port map (
            O => \N__35090\,
            I => \N__35079\
        );

    \I__6790\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35079\
        );

    \I__6789\ : Odrv4
    port map (
            O => \N__35086\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__35079\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__6787\ : InMux
    port map (
            O => \N__35074\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__6786\ : CascadeMux
    port map (
            O => \N__35071\,
            I => \N__35067\
        );

    \I__6785\ : CascadeMux
    port map (
            O => \N__35070\,
            I => \N__35064\
        );

    \I__6784\ : InMux
    port map (
            O => \N__35067\,
            I => \N__35059\
        );

    \I__6783\ : InMux
    port map (
            O => \N__35064\,
            I => \N__35059\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__35059\,
            I => \N__35055\
        );

    \I__6781\ : InMux
    port map (
            O => \N__35058\,
            I => \N__35052\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__35055\,
            I => \N__35049\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__35052\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__6778\ : Odrv4
    port map (
            O => \N__35049\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__6777\ : InMux
    port map (
            O => \N__35044\,
            I => \N__35041\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__35041\,
            I => \N__35035\
        );

    \I__6775\ : InMux
    port map (
            O => \N__35040\,
            I => \N__35032\
        );

    \I__6774\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35029\
        );

    \I__6773\ : InMux
    port map (
            O => \N__35038\,
            I => \N__35026\
        );

    \I__6772\ : Odrv4
    port map (
            O => \N__35035\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__35032\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__35029\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__35026\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__6768\ : InMux
    port map (
            O => \N__35017\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__6767\ : CascadeMux
    port map (
            O => \N__35014\,
            I => \N__35010\
        );

    \I__6766\ : InMux
    port map (
            O => \N__35013\,
            I => \N__35007\
        );

    \I__6765\ : InMux
    port map (
            O => \N__35010\,
            I => \N__35004\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__35007\,
            I => \N__34998\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__35004\,
            I => \N__34998\
        );

    \I__6762\ : InMux
    port map (
            O => \N__35003\,
            I => \N__34995\
        );

    \I__6761\ : Span4Mux_v
    port map (
            O => \N__34998\,
            I => \N__34992\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__34995\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__6759\ : Odrv4
    port map (
            O => \N__34992\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__34987\,
            I => \N__34983\
        );

    \I__6757\ : CascadeMux
    port map (
            O => \N__34986\,
            I => \N__34979\
        );

    \I__6756\ : InMux
    port map (
            O => \N__34983\,
            I => \N__34976\
        );

    \I__6755\ : CascadeMux
    port map (
            O => \N__34982\,
            I => \N__34973\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34979\,
            I => \N__34969\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__34976\,
            I => \N__34966\
        );

    \I__6752\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34963\
        );

    \I__6751\ : InMux
    port map (
            O => \N__34972\,
            I => \N__34960\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__34969\,
            I => \N__34957\
        );

    \I__6749\ : Odrv4
    port map (
            O => \N__34966\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__34963\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__34960\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__6746\ : Odrv4
    port map (
            O => \N__34957\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__6745\ : InMux
    port map (
            O => \N__34948\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__6744\ : InMux
    port map (
            O => \N__34945\,
            I => \N__34939\
        );

    \I__6743\ : InMux
    port map (
            O => \N__34944\,
            I => \N__34939\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__34939\,
            I => \N__34935\
        );

    \I__6741\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34932\
        );

    \I__6740\ : Span4Mux_v
    port map (
            O => \N__34935\,
            I => \N__34929\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__34932\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__6738\ : Odrv4
    port map (
            O => \N__34929\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__6737\ : InMux
    port map (
            O => \N__34924\,
            I => \N__34921\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__34921\,
            I => \N__34917\
        );

    \I__6735\ : CascadeMux
    port map (
            O => \N__34920\,
            I => \N__34913\
        );

    \I__6734\ : Span4Mux_h
    port map (
            O => \N__34917\,
            I => \N__34909\
        );

    \I__6733\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34906\
        );

    \I__6732\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34901\
        );

    \I__6731\ : InMux
    port map (
            O => \N__34912\,
            I => \N__34901\
        );

    \I__6730\ : Odrv4
    port map (
            O => \N__34909\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__34906\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__34901\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__6727\ : InMux
    port map (
            O => \N__34894\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__6726\ : InMux
    port map (
            O => \N__34891\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__6725\ : InMux
    port map (
            O => \N__34888\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__6724\ : InMux
    port map (
            O => \N__34885\,
            I => \bfn_14_24_0_\
        );

    \I__6723\ : InMux
    port map (
            O => \N__34882\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__6722\ : InMux
    port map (
            O => \N__34879\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__6721\ : InMux
    port map (
            O => \N__34876\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__6720\ : InMux
    port map (
            O => \N__34873\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__6719\ : InMux
    port map (
            O => \N__34870\,
            I => \N__34840\
        );

    \I__6718\ : InMux
    port map (
            O => \N__34869\,
            I => \N__34840\
        );

    \I__6717\ : InMux
    port map (
            O => \N__34868\,
            I => \N__34840\
        );

    \I__6716\ : InMux
    port map (
            O => \N__34867\,
            I => \N__34840\
        );

    \I__6715\ : InMux
    port map (
            O => \N__34866\,
            I => \N__34831\
        );

    \I__6714\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34831\
        );

    \I__6713\ : InMux
    port map (
            O => \N__34864\,
            I => \N__34831\
        );

    \I__6712\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34831\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34862\,
            I => \N__34826\
        );

    \I__6710\ : InMux
    port map (
            O => \N__34861\,
            I => \N__34826\
        );

    \I__6709\ : InMux
    port map (
            O => \N__34860\,
            I => \N__34809\
        );

    \I__6708\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34809\
        );

    \I__6707\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34809\
        );

    \I__6706\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34809\
        );

    \I__6705\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34800\
        );

    \I__6704\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34800\
        );

    \I__6703\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34800\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34853\,
            I => \N__34800\
        );

    \I__6701\ : InMux
    port map (
            O => \N__34852\,
            I => \N__34791\
        );

    \I__6700\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34791\
        );

    \I__6699\ : InMux
    port map (
            O => \N__34850\,
            I => \N__34791\
        );

    \I__6698\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34791\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__34840\,
            I => \N__34784\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__34831\,
            I => \N__34784\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__34826\,
            I => \N__34784\
        );

    \I__6694\ : InMux
    port map (
            O => \N__34825\,
            I => \N__34775\
        );

    \I__6693\ : InMux
    port map (
            O => \N__34824\,
            I => \N__34775\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34823\,
            I => \N__34775\
        );

    \I__6691\ : InMux
    port map (
            O => \N__34822\,
            I => \N__34775\
        );

    \I__6690\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34766\
        );

    \I__6689\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34766\
        );

    \I__6688\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34766\
        );

    \I__6687\ : InMux
    port map (
            O => \N__34818\,
            I => \N__34766\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__34809\,
            I => \N__34759\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__34800\,
            I => \N__34759\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__34791\,
            I => \N__34759\
        );

    \I__6683\ : Span4Mux_v
    port map (
            O => \N__34784\,
            I => \N__34756\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__34775\,
            I => \N__34747\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__34766\,
            I => \N__34747\
        );

    \I__6680\ : Span4Mux_v
    port map (
            O => \N__34759\,
            I => \N__34747\
        );

    \I__6679\ : Span4Mux_h
    port map (
            O => \N__34756\,
            I => \N__34747\
        );

    \I__6678\ : Odrv4
    port map (
            O => \N__34747\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__6677\ : InMux
    port map (
            O => \N__34744\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__6676\ : CEMux
    port map (
            O => \N__34741\,
            I => \N__34736\
        );

    \I__6675\ : CEMux
    port map (
            O => \N__34740\,
            I => \N__34733\
        );

    \I__6674\ : CEMux
    port map (
            O => \N__34739\,
            I => \N__34730\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__34736\,
            I => \N__34727\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__34733\,
            I => \N__34721\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__34730\,
            I => \N__34721\
        );

    \I__6670\ : Span4Mux_v
    port map (
            O => \N__34727\,
            I => \N__34718\
        );

    \I__6669\ : CEMux
    port map (
            O => \N__34726\,
            I => \N__34715\
        );

    \I__6668\ : Span4Mux_v
    port map (
            O => \N__34721\,
            I => \N__34712\
        );

    \I__6667\ : Span4Mux_h
    port map (
            O => \N__34718\,
            I => \N__34707\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__34715\,
            I => \N__34707\
        );

    \I__6665\ : Span4Mux_h
    port map (
            O => \N__34712\,
            I => \N__34702\
        );

    \I__6664\ : Span4Mux_h
    port map (
            O => \N__34707\,
            I => \N__34702\
        );

    \I__6663\ : Span4Mux_v
    port map (
            O => \N__34702\,
            I => \N__34699\
        );

    \I__6662\ : Span4Mux_v
    port map (
            O => \N__34699\,
            I => \N__34696\
        );

    \I__6661\ : Odrv4
    port map (
            O => \N__34696\,
            I => \delay_measurement_inst.delay_hc_timer.N_303_i\
        );

    \I__6660\ : InMux
    port map (
            O => \N__34693\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__6659\ : InMux
    port map (
            O => \N__34690\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34687\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__6657\ : InMux
    port map (
            O => \N__34684\,
            I => \bfn_14_23_0_\
        );

    \I__6656\ : InMux
    port map (
            O => \N__34681\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__6655\ : InMux
    port map (
            O => \N__34678\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__6654\ : InMux
    port map (
            O => \N__34675\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__6653\ : InMux
    port map (
            O => \N__34672\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__6652\ : InMux
    port map (
            O => \N__34669\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__6651\ : InMux
    port map (
            O => \N__34666\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__6650\ : InMux
    port map (
            O => \N__34663\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__6649\ : InMux
    port map (
            O => \N__34660\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__6648\ : InMux
    port map (
            O => \N__34657\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__6647\ : InMux
    port map (
            O => \N__34654\,
            I => \bfn_14_22_0_\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34651\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__6645\ : InMux
    port map (
            O => \N__34648\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__6644\ : InMux
    port map (
            O => \N__34645\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__6643\ : InMux
    port map (
            O => \N__34642\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__6642\ : InMux
    port map (
            O => \N__34639\,
            I => \N__34636\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__34636\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__6640\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34630\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__34630\,
            I => \N__34627\
        );

    \I__6638\ : Odrv4
    port map (
            O => \N__34627\,
            I => \current_shift_inst.control_input_1_axb_19\
        );

    \I__6637\ : InMux
    port map (
            O => \N__34624\,
            I => \N__34621\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__34621\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__6635\ : InMux
    port map (
            O => \N__34618\,
            I => \N__34615\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__34615\,
            I => \current_shift_inst.control_input_1_axb_24\
        );

    \I__6633\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34609\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__34609\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__6631\ : InMux
    port map (
            O => \N__34606\,
            I => \N__34603\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__34603\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__6629\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34597\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__34597\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__6627\ : InMux
    port map (
            O => \N__34594\,
            I => \bfn_14_21_0_\
        );

    \I__6626\ : InMux
    port map (
            O => \N__34591\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__6625\ : InMux
    port map (
            O => \N__34588\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__6624\ : InMux
    port map (
            O => \N__34585\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__6623\ : InMux
    port map (
            O => \N__34582\,
            I => \N__34579\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__34579\,
            I => \N__34576\
        );

    \I__6621\ : Odrv4
    port map (
            O => \N__34576\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__6620\ : InMux
    port map (
            O => \N__34573\,
            I => \N__34570\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__34570\,
            I => \current_shift_inst.control_input_1_axb_16\
        );

    \I__6618\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34564\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__34564\,
            I => \N__34561\
        );

    \I__6616\ : Span4Mux_h
    port map (
            O => \N__34561\,
            I => \N__34558\
        );

    \I__6615\ : Odrv4
    port map (
            O => \N__34558\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__6614\ : InMux
    port map (
            O => \N__34555\,
            I => \N__34552\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__34552\,
            I => \current_shift_inst.control_input_1_axb_23\
        );

    \I__6612\ : InMux
    port map (
            O => \N__34549\,
            I => \N__34546\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__34546\,
            I => \N__34543\
        );

    \I__6610\ : Odrv4
    port map (
            O => \N__34543\,
            I => \current_shift_inst.un38_control_input_0_s0_7\
        );

    \I__6609\ : InMux
    port map (
            O => \N__34540\,
            I => \N__34537\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__34537\,
            I => \N__34534\
        );

    \I__6607\ : Odrv12
    port map (
            O => \N__34534\,
            I => \current_shift_inst.control_input_1_axb_1\
        );

    \I__6606\ : InMux
    port map (
            O => \N__34531\,
            I => \N__34528\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__34528\,
            I => \N__34525\
        );

    \I__6604\ : Odrv4
    port map (
            O => \N__34525\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__6603\ : InMux
    port map (
            O => \N__34522\,
            I => \N__34519\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__34519\,
            I => \N__34516\
        );

    \I__6601\ : Odrv4
    port map (
            O => \N__34516\,
            I => \current_shift_inst.control_input_1_axb_21\
        );

    \I__6600\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34510\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__34510\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\
        );

    \I__6598\ : CascadeMux
    port map (
            O => \N__34507\,
            I => \N__34504\
        );

    \I__6597\ : InMux
    port map (
            O => \N__34504\,
            I => \N__34501\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__34501\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\
        );

    \I__6595\ : InMux
    port map (
            O => \N__34498\,
            I => \N__34495\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__34495\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__6593\ : InMux
    port map (
            O => \N__34492\,
            I => \N__34489\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__34489\,
            I => \N__34486\
        );

    \I__6591\ : Odrv4
    port map (
            O => \N__34486\,
            I => \current_shift_inst.control_input_1_axb_18\
        );

    \I__6590\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34480\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__34480\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__6588\ : InMux
    port map (
            O => \N__34477\,
            I => \N__34474\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__34474\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__6586\ : InMux
    port map (
            O => \N__34471\,
            I => \N__34468\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__34468\,
            I => \N__34465\
        );

    \I__6584\ : Odrv4
    port map (
            O => \N__34465\,
            I => \current_shift_inst.control_input_1_axb_20\
        );

    \I__6583\ : InMux
    port map (
            O => \N__34462\,
            I => \N__34459\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__34459\,
            I => \N__34456\
        );

    \I__6581\ : Span4Mux_v
    port map (
            O => \N__34456\,
            I => \N__34453\
        );

    \I__6580\ : Span4Mux_h
    port map (
            O => \N__34453\,
            I => \N__34450\
        );

    \I__6579\ : Odrv4
    port map (
            O => \N__34450\,
            I => \current_shift_inst.control_inputZ0Z_21\
        );

    \I__6578\ : InMux
    port map (
            O => \N__34447\,
            I => \current_shift_inst.control_input_1_cry_20\
        );

    \I__6577\ : InMux
    port map (
            O => \N__34444\,
            I => \N__34441\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__34441\,
            I => \N__34438\
        );

    \I__6575\ : Span4Mux_h
    port map (
            O => \N__34438\,
            I => \N__34435\
        );

    \I__6574\ : Odrv4
    port map (
            O => \N__34435\,
            I => \current_shift_inst.control_inputZ0Z_22\
        );

    \I__6573\ : InMux
    port map (
            O => \N__34432\,
            I => \current_shift_inst.control_input_1_cry_21\
        );

    \I__6572\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34426\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__34426\,
            I => \N__34423\
        );

    \I__6570\ : Odrv12
    port map (
            O => \N__34423\,
            I => \current_shift_inst.control_inputZ0Z_23\
        );

    \I__6569\ : InMux
    port map (
            O => \N__34420\,
            I => \current_shift_inst.control_input_1_cry_22\
        );

    \I__6568\ : InMux
    port map (
            O => \N__34417\,
            I => \N__34414\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__34414\,
            I => \N__34411\
        );

    \I__6566\ : Span4Mux_v
    port map (
            O => \N__34411\,
            I => \N__34408\
        );

    \I__6565\ : Odrv4
    port map (
            O => \N__34408\,
            I => \current_shift_inst.control_inputZ0Z_24\
        );

    \I__6564\ : InMux
    port map (
            O => \N__34405\,
            I => \bfn_14_18_0_\
        );

    \I__6563\ : InMux
    port map (
            O => \N__34402\,
            I => \N__34399\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__34399\,
            I => \N__34396\
        );

    \I__6561\ : Span4Mux_h
    port map (
            O => \N__34396\,
            I => \N__34393\
        );

    \I__6560\ : Odrv4
    port map (
            O => \N__34393\,
            I => \current_shift_inst.control_input_1_axb_25\
        );

    \I__6559\ : InMux
    port map (
            O => \N__34390\,
            I => \current_shift_inst.control_input_1_cry_24\
        );

    \I__6558\ : InMux
    port map (
            O => \N__34387\,
            I => \N__34381\
        );

    \I__6557\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34381\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__34381\,
            I => \N__34378\
        );

    \I__6555\ : Span4Mux_v
    port map (
            O => \N__34378\,
            I => \N__34375\
        );

    \I__6554\ : Odrv4
    port map (
            O => \N__34375\,
            I => \current_shift_inst.control_inputZ0Z_25\
        );

    \I__6553\ : InMux
    port map (
            O => \N__34372\,
            I => \N__34369\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__34369\,
            I => \N__34366\
        );

    \I__6551\ : Odrv4
    port map (
            O => \N__34366\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__6550\ : InMux
    port map (
            O => \N__34363\,
            I => \N__34360\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__34360\,
            I => \current_shift_inst.control_input_1_axb_22\
        );

    \I__6548\ : CascadeMux
    port map (
            O => \N__34357\,
            I => \N__34353\
        );

    \I__6547\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34350\
        );

    \I__6546\ : InMux
    port map (
            O => \N__34353\,
            I => \N__34347\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__34350\,
            I => \N__34342\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__34347\,
            I => \N__34342\
        );

    \I__6543\ : Odrv4
    port map (
            O => \N__34342\,
            I => \current_shift_inst.N_1355_i\
        );

    \I__6542\ : InMux
    port map (
            O => \N__34339\,
            I => \N__34336\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__34336\,
            I => \current_shift_inst.un38_control_input_0_s0_6\
        );

    \I__6540\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34330\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__34330\,
            I => \N__34327\
        );

    \I__6538\ : Odrv4
    port map (
            O => \N__34327\,
            I => \current_shift_inst.control_input_1_axb_0\
        );

    \I__6537\ : InMux
    port map (
            O => \N__34324\,
            I => \N__34321\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__34321\,
            I => \N__34318\
        );

    \I__6535\ : Odrv4
    port map (
            O => \N__34318\,
            I => \current_shift_inst.control_input_1_axb_13\
        );

    \I__6534\ : InMux
    port map (
            O => \N__34315\,
            I => \N__34312\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__34312\,
            I => \N__34309\
        );

    \I__6532\ : Odrv12
    port map (
            O => \N__34309\,
            I => \current_shift_inst.control_inputZ0Z_13\
        );

    \I__6531\ : InMux
    port map (
            O => \N__34306\,
            I => \current_shift_inst.control_input_1_cry_12\
        );

    \I__6530\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34300\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__34300\,
            I => \current_shift_inst.control_input_1_axb_14\
        );

    \I__6528\ : InMux
    port map (
            O => \N__34297\,
            I => \N__34294\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__34294\,
            I => \N__34291\
        );

    \I__6526\ : Odrv12
    port map (
            O => \N__34291\,
            I => \current_shift_inst.control_inputZ0Z_14\
        );

    \I__6525\ : InMux
    port map (
            O => \N__34288\,
            I => \current_shift_inst.control_input_1_cry_13\
        );

    \I__6524\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34282\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__34282\,
            I => \current_shift_inst.control_input_1_axb_15\
        );

    \I__6522\ : InMux
    port map (
            O => \N__34279\,
            I => \N__34276\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__34276\,
            I => \N__34273\
        );

    \I__6520\ : Odrv12
    port map (
            O => \N__34273\,
            I => \current_shift_inst.control_inputZ0Z_15\
        );

    \I__6519\ : InMux
    port map (
            O => \N__34270\,
            I => \current_shift_inst.control_input_1_cry_14\
        );

    \I__6518\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34264\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__34264\,
            I => \N__34261\
        );

    \I__6516\ : Odrv12
    port map (
            O => \N__34261\,
            I => \current_shift_inst.control_inputZ0Z_16\
        );

    \I__6515\ : InMux
    port map (
            O => \N__34258\,
            I => \bfn_14_17_0_\
        );

    \I__6514\ : InMux
    port map (
            O => \N__34255\,
            I => \N__34252\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__34252\,
            I => \current_shift_inst.control_input_1_axb_17\
        );

    \I__6512\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34246\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__34246\,
            I => \N__34243\
        );

    \I__6510\ : Span12Mux_v
    port map (
            O => \N__34243\,
            I => \N__34240\
        );

    \I__6509\ : Odrv12
    port map (
            O => \N__34240\,
            I => \current_shift_inst.control_inputZ0Z_17\
        );

    \I__6508\ : InMux
    port map (
            O => \N__34237\,
            I => \current_shift_inst.control_input_1_cry_16\
        );

    \I__6507\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34231\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__34231\,
            I => \N__34228\
        );

    \I__6505\ : Odrv12
    port map (
            O => \N__34228\,
            I => \current_shift_inst.control_inputZ0Z_18\
        );

    \I__6504\ : InMux
    port map (
            O => \N__34225\,
            I => \current_shift_inst.control_input_1_cry_17\
        );

    \I__6503\ : InMux
    port map (
            O => \N__34222\,
            I => \N__34219\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__34219\,
            I => \N__34216\
        );

    \I__6501\ : Odrv12
    port map (
            O => \N__34216\,
            I => \current_shift_inst.control_inputZ0Z_19\
        );

    \I__6500\ : InMux
    port map (
            O => \N__34213\,
            I => \current_shift_inst.control_input_1_cry_18\
        );

    \I__6499\ : InMux
    port map (
            O => \N__34210\,
            I => \N__34207\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__34207\,
            I => \N__34204\
        );

    \I__6497\ : Odrv12
    port map (
            O => \N__34204\,
            I => \current_shift_inst.control_inputZ0Z_20\
        );

    \I__6496\ : InMux
    port map (
            O => \N__34201\,
            I => \current_shift_inst.control_input_1_cry_19\
        );

    \I__6495\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34195\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__34195\,
            I => \N__34192\
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__34192\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__6492\ : InMux
    port map (
            O => \N__34189\,
            I => \current_shift_inst.control_input_1_cry_4\
        );

    \I__6491\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34183\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__34183\,
            I => \current_shift_inst.control_input_1_axb_6\
        );

    \I__6489\ : InMux
    port map (
            O => \N__34180\,
            I => \N__34177\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__34177\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__6487\ : InMux
    port map (
            O => \N__34174\,
            I => \current_shift_inst.control_input_1_cry_5\
        );

    \I__6486\ : InMux
    port map (
            O => \N__34171\,
            I => \N__34168\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__34168\,
            I => \N__34165\
        );

    \I__6484\ : Odrv12
    port map (
            O => \N__34165\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__6483\ : InMux
    port map (
            O => \N__34162\,
            I => \current_shift_inst.control_input_1_cry_6\
        );

    \I__6482\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34156\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__34156\,
            I => \current_shift_inst.control_input_1_axb_8\
        );

    \I__6480\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34150\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__34150\,
            I => \N__34147\
        );

    \I__6478\ : Odrv12
    port map (
            O => \N__34147\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__6477\ : InMux
    port map (
            O => \N__34144\,
            I => \bfn_14_16_0_\
        );

    \I__6476\ : InMux
    port map (
            O => \N__34141\,
            I => \N__34138\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__34138\,
            I => \current_shift_inst.control_input_1_axb_9\
        );

    \I__6474\ : InMux
    port map (
            O => \N__34135\,
            I => \N__34132\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__34132\,
            I => \N__34129\
        );

    \I__6472\ : Span4Mux_h
    port map (
            O => \N__34129\,
            I => \N__34126\
        );

    \I__6471\ : Span4Mux_v
    port map (
            O => \N__34126\,
            I => \N__34123\
        );

    \I__6470\ : Odrv4
    port map (
            O => \N__34123\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__6469\ : InMux
    port map (
            O => \N__34120\,
            I => \current_shift_inst.control_input_1_cry_8\
        );

    \I__6468\ : InMux
    port map (
            O => \N__34117\,
            I => \N__34114\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__34114\,
            I => \N__34111\
        );

    \I__6466\ : Odrv4
    port map (
            O => \N__34111\,
            I => \current_shift_inst.control_input_1_axb_10\
        );

    \I__6465\ : InMux
    port map (
            O => \N__34108\,
            I => \N__34105\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__34105\,
            I => \N__34102\
        );

    \I__6463\ : Odrv12
    port map (
            O => \N__34102\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__6462\ : InMux
    port map (
            O => \N__34099\,
            I => \current_shift_inst.control_input_1_cry_9\
        );

    \I__6461\ : InMux
    port map (
            O => \N__34096\,
            I => \N__34093\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__34093\,
            I => \current_shift_inst.control_input_1_axb_11\
        );

    \I__6459\ : InMux
    port map (
            O => \N__34090\,
            I => \N__34087\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__34087\,
            I => \N__34084\
        );

    \I__6457\ : Odrv12
    port map (
            O => \N__34084\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__6456\ : InMux
    port map (
            O => \N__34081\,
            I => \current_shift_inst.control_input_1_cry_10\
        );

    \I__6455\ : InMux
    port map (
            O => \N__34078\,
            I => \N__34075\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__34075\,
            I => \current_shift_inst.control_input_1_axb_12\
        );

    \I__6453\ : InMux
    port map (
            O => \N__34072\,
            I => \N__34069\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__34069\,
            I => \N__34066\
        );

    \I__6451\ : Odrv4
    port map (
            O => \N__34066\,
            I => \current_shift_inst.control_inputZ0Z_12\
        );

    \I__6450\ : InMux
    port map (
            O => \N__34063\,
            I => \current_shift_inst.control_input_1_cry_11\
        );

    \I__6449\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34057\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__34057\,
            I => \N__34054\
        );

    \I__6447\ : Span4Mux_h
    port map (
            O => \N__34054\,
            I => \N__34051\
        );

    \I__6446\ : Odrv4
    port map (
            O => \N__34051\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\
        );

    \I__6445\ : InMux
    port map (
            O => \N__34048\,
            I => \N__34035\
        );

    \I__6444\ : InMux
    port map (
            O => \N__34047\,
            I => \N__34035\
        );

    \I__6443\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34035\
        );

    \I__6442\ : InMux
    port map (
            O => \N__34045\,
            I => \N__34030\
        );

    \I__6441\ : InMux
    port map (
            O => \N__34044\,
            I => \N__34030\
        );

    \I__6440\ : CascadeMux
    port map (
            O => \N__34043\,
            I => \N__34027\
        );

    \I__6439\ : InMux
    port map (
            O => \N__34042\,
            I => \N__34022\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__34035\,
            I => \N__34016\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__34030\,
            I => \N__34016\
        );

    \I__6436\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34013\
        );

    \I__6435\ : InMux
    port map (
            O => \N__34026\,
            I => \N__34010\
        );

    \I__6434\ : InMux
    port map (
            O => \N__34025\,
            I => \N__34007\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__34022\,
            I => \N__34004\
        );

    \I__6432\ : InMux
    port map (
            O => \N__34021\,
            I => \N__34001\
        );

    \I__6431\ : Span4Mux_h
    port map (
            O => \N__34016\,
            I => \N__33996\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__34013\,
            I => \N__33996\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__34010\,
            I => measured_delay_tr_15
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__34007\,
            I => measured_delay_tr_15
        );

    \I__6427\ : Odrv4
    port map (
            O => \N__34004\,
            I => measured_delay_tr_15
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__34001\,
            I => measured_delay_tr_15
        );

    \I__6425\ : Odrv4
    port map (
            O => \N__33996\,
            I => measured_delay_tr_15
        );

    \I__6424\ : InMux
    port map (
            O => \N__33985\,
            I => \N__33980\
        );

    \I__6423\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33975\
        );

    \I__6422\ : InMux
    port map (
            O => \N__33983\,
            I => \N__33975\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__33980\,
            I => \N__33972\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__33975\,
            I => \N__33969\
        );

    \I__6419\ : Span4Mux_h
    port map (
            O => \N__33972\,
            I => \N__33963\
        );

    \I__6418\ : Span4Mux_h
    port map (
            O => \N__33969\,
            I => \N__33960\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33957\
        );

    \I__6416\ : InMux
    port map (
            O => \N__33967\,
            I => \N__33952\
        );

    \I__6415\ : InMux
    port map (
            O => \N__33966\,
            I => \N__33952\
        );

    \I__6414\ : Odrv4
    port map (
            O => \N__33963\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__6413\ : Odrv4
    port map (
            O => \N__33960\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__33957\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__33952\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__6410\ : CascadeMux
    port map (
            O => \N__33943\,
            I => \N__33940\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33937\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__33937\,
            I => \N__33934\
        );

    \I__6407\ : Span4Mux_h
    port map (
            O => \N__33934\,
            I => \N__33931\
        );

    \I__6406\ : Odrv4
    port map (
            O => \N__33931\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__6405\ : CEMux
    port map (
            O => \N__33928\,
            I => \N__33922\
        );

    \I__6404\ : CEMux
    port map (
            O => \N__33927\,
            I => \N__33918\
        );

    \I__6403\ : CEMux
    port map (
            O => \N__33926\,
            I => \N__33914\
        );

    \I__6402\ : CEMux
    port map (
            O => \N__33925\,
            I => \N__33911\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__33922\,
            I => \N__33908\
        );

    \I__6400\ : CEMux
    port map (
            O => \N__33921\,
            I => \N__33905\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__33918\,
            I => \N__33902\
        );

    \I__6398\ : CEMux
    port map (
            O => \N__33917\,
            I => \N__33899\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__33914\,
            I => \N__33896\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__33911\,
            I => \N__33893\
        );

    \I__6395\ : Span4Mux_v
    port map (
            O => \N__33908\,
            I => \N__33890\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__33905\,
            I => \N__33887\
        );

    \I__6393\ : Span4Mux_h
    port map (
            O => \N__33902\,
            I => \N__33884\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33879\
        );

    \I__6391\ : Span4Mux_h
    port map (
            O => \N__33896\,
            I => \N__33879\
        );

    \I__6390\ : Span4Mux_h
    port map (
            O => \N__33893\,
            I => \N__33876\
        );

    \I__6389\ : Span4Mux_h
    port map (
            O => \N__33890\,
            I => \N__33871\
        );

    \I__6388\ : Span4Mux_h
    port map (
            O => \N__33887\,
            I => \N__33871\
        );

    \I__6387\ : Odrv4
    port map (
            O => \N__33884\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__6386\ : Odrv4
    port map (
            O => \N__33879\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__33876\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__6384\ : Odrv4
    port map (
            O => \N__33871\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__6383\ : InMux
    port map (
            O => \N__33862\,
            I => \N__33859\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__33859\,
            I => \N__33856\
        );

    \I__6381\ : Span4Mux_h
    port map (
            O => \N__33856\,
            I => \N__33853\
        );

    \I__6380\ : Odrv4
    port map (
            O => \N__33853\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__6379\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33847\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__33847\,
            I => \N__33844\
        );

    \I__6377\ : Span4Mux_h
    port map (
            O => \N__33844\,
            I => \N__33841\
        );

    \I__6376\ : Odrv4
    port map (
            O => \N__33841\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\
        );

    \I__6375\ : InMux
    port map (
            O => \N__33838\,
            I => \N__33835\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__33835\,
            I => \N__33831\
        );

    \I__6373\ : InMux
    port map (
            O => \N__33834\,
            I => \N__33828\
        );

    \I__6372\ : Span4Mux_v
    port map (
            O => \N__33831\,
            I => \N__33823\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__33828\,
            I => \N__33823\
        );

    \I__6370\ : Span4Mux_v
    port map (
            O => \N__33823\,
            I => \N__33820\
        );

    \I__6369\ : Odrv4
    port map (
            O => \N__33820\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__6368\ : InMux
    port map (
            O => \N__33817\,
            I => \N__33814\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__33814\,
            I => \N__33811\
        );

    \I__6366\ : Odrv4
    port map (
            O => \N__33811\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__6365\ : InMux
    port map (
            O => \N__33808\,
            I => \current_shift_inst.control_input_1_cry_0\
        );

    \I__6364\ : InMux
    port map (
            O => \N__33805\,
            I => \N__33802\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__33802\,
            I => \current_shift_inst.control_input_1_axb_2\
        );

    \I__6362\ : InMux
    port map (
            O => \N__33799\,
            I => \N__33796\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__33796\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__6360\ : InMux
    port map (
            O => \N__33793\,
            I => \current_shift_inst.control_input_1_cry_1\
        );

    \I__6359\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33787\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__33787\,
            I => \current_shift_inst.control_input_1_axb_3\
        );

    \I__6357\ : InMux
    port map (
            O => \N__33784\,
            I => \N__33781\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__33781\,
            I => \N__33778\
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__33778\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__6354\ : InMux
    port map (
            O => \N__33775\,
            I => \current_shift_inst.control_input_1_cry_2\
        );

    \I__6353\ : InMux
    port map (
            O => \N__33772\,
            I => \N__33769\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__33769\,
            I => \current_shift_inst.control_input_1_axb_4\
        );

    \I__6351\ : InMux
    port map (
            O => \N__33766\,
            I => \N__33763\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__33763\,
            I => \N__33760\
        );

    \I__6349\ : Span4Mux_v
    port map (
            O => \N__33760\,
            I => \N__33757\
        );

    \I__6348\ : Span4Mux_h
    port map (
            O => \N__33757\,
            I => \N__33754\
        );

    \I__6347\ : Odrv4
    port map (
            O => \N__33754\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__6346\ : InMux
    port map (
            O => \N__33751\,
            I => \current_shift_inst.control_input_1_cry_3\
        );

    \I__6345\ : InMux
    port map (
            O => \N__33748\,
            I => \N__33745\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__33745\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__6343\ : InMux
    port map (
            O => \N__33742\,
            I => \N__33739\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__33739\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__6341\ : CascadeMux
    port map (
            O => \N__33736\,
            I => \N__33733\
        );

    \I__6340\ : InMux
    port map (
            O => \N__33733\,
            I => \N__33730\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__33730\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\
        );

    \I__6338\ : CascadeMux
    port map (
            O => \N__33727\,
            I => \N__33724\
        );

    \I__6337\ : InMux
    port map (
            O => \N__33724\,
            I => \N__33721\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__33721\,
            I => \N__33718\
        );

    \I__6335\ : Odrv4
    port map (
            O => \N__33718\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__6334\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33712\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__33712\,
            I => \N__33709\
        );

    \I__6332\ : Odrv4
    port map (
            O => \N__33709\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\
        );

    \I__6331\ : InMux
    port map (
            O => \N__33706\,
            I => \N__33703\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__33703\,
            I => \N__33700\
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__33700\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__6328\ : InMux
    port map (
            O => \N__33697\,
            I => \N__33694\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__33694\,
            I => \N__33691\
        );

    \I__6326\ : Odrv4
    port map (
            O => \N__33691\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__6325\ : InMux
    port map (
            O => \N__33688\,
            I => \N__33685\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__33685\,
            I => \N__33682\
        );

    \I__6323\ : Span4Mux_h
    port map (
            O => \N__33682\,
            I => \N__33679\
        );

    \I__6322\ : Odrv4
    port map (
            O => \N__33679\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\
        );

    \I__6321\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33673\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__33673\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\
        );

    \I__6319\ : InMux
    port map (
            O => \N__33670\,
            I => \N__33667\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__33667\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__6317\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33661\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__33661\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__6315\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33655\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__33655\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\
        );

    \I__6313\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33649\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__33649\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__6311\ : InMux
    port map (
            O => \N__33646\,
            I => \N__33643\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__33643\,
            I => \N__33640\
        );

    \I__6309\ : Odrv12
    port map (
            O => \N__33640\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__6308\ : InMux
    port map (
            O => \N__33637\,
            I => \N__33634\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__33634\,
            I => \N__33631\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__33631\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__6305\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33625\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__33625\,
            I => \N__33622\
        );

    \I__6303\ : Odrv4
    port map (
            O => \N__33622\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__6302\ : InMux
    port map (
            O => \N__33619\,
            I => \N__33616\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__33616\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\
        );

    \I__6300\ : InMux
    port map (
            O => \N__33613\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\
        );

    \I__6299\ : InMux
    port map (
            O => \N__33610\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\
        );

    \I__6298\ : InMux
    port map (
            O => \N__33607\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\
        );

    \I__6297\ : InMux
    port map (
            O => \N__33604\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_31\
        );

    \I__6296\ : InMux
    port map (
            O => \N__33601\,
            I => \N__33598\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__33598\,
            I => \N__33595\
        );

    \I__6294\ : Odrv4
    port map (
            O => \N__33595\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__6293\ : InMux
    port map (
            O => \N__33592\,
            I => \N__33589\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__33589\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__6291\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33583\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__33583\,
            I => \N__33580\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__33580\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__6288\ : InMux
    port map (
            O => \N__33577\,
            I => \N__33574\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__33574\,
            I => \N__33571\
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__33571\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__6285\ : InMux
    port map (
            O => \N__33568\,
            I => \N__33565\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__33565\,
            I => \N__33562\
        );

    \I__6283\ : Odrv4
    port map (
            O => \N__33562\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__6282\ : InMux
    port map (
            O => \N__33559\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\
        );

    \I__6281\ : InMux
    port map (
            O => \N__33556\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\
        );

    \I__6280\ : InMux
    port map (
            O => \N__33553\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\
        );

    \I__6279\ : InMux
    port map (
            O => \N__33550\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\
        );

    \I__6278\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33544\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__33544\,
            I => \N__33541\
        );

    \I__6276\ : Span4Mux_h
    port map (
            O => \N__33541\,
            I => \N__33538\
        );

    \I__6275\ : Odrv4
    port map (
            O => \N__33538\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__6274\ : InMux
    port map (
            O => \N__33535\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\
        );

    \I__6273\ : InMux
    port map (
            O => \N__33532\,
            I => \bfn_14_10_0_\
        );

    \I__6272\ : InMux
    port map (
            O => \N__33529\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\
        );

    \I__6271\ : InMux
    port map (
            O => \N__33526\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\
        );

    \I__6270\ : InMux
    port map (
            O => \N__33523\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\
        );

    \I__6269\ : InMux
    port map (
            O => \N__33520\,
            I => \N__33517\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__33517\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\
        );

    \I__6267\ : InMux
    port map (
            O => \N__33514\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\
        );

    \I__6266\ : InMux
    port map (
            O => \N__33511\,
            I => \N__33508\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__33508\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\
        );

    \I__6264\ : InMux
    port map (
            O => \N__33505\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\
        );

    \I__6263\ : InMux
    port map (
            O => \N__33502\,
            I => \N__33499\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__33499\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__6261\ : InMux
    port map (
            O => \N__33496\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\
        );

    \I__6260\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33490\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__33490\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__6258\ : InMux
    port map (
            O => \N__33487\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\
        );

    \I__6257\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33481\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__33481\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__6255\ : InMux
    port map (
            O => \N__33478\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\
        );

    \I__6254\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33472\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__33472\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33469\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\
        );

    \I__6251\ : InMux
    port map (
            O => \N__33466\,
            I => \N__33463\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__33463\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__6249\ : InMux
    port map (
            O => \N__33460\,
            I => \bfn_14_9_0_\
        );

    \I__6248\ : InMux
    port map (
            O => \N__33457\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\
        );

    \I__6247\ : InMux
    port map (
            O => \N__33454\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\
        );

    \I__6246\ : InMux
    port map (
            O => \N__33451\,
            I => \N__33447\
        );

    \I__6245\ : InMux
    port map (
            O => \N__33450\,
            I => \N__33444\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__33447\,
            I => \N__33441\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__33444\,
            I => \N__33438\
        );

    \I__6242\ : Span4Mux_v
    port map (
            O => \N__33441\,
            I => \N__33435\
        );

    \I__6241\ : Span4Mux_h
    port map (
            O => \N__33438\,
            I => \N__33432\
        );

    \I__6240\ : Odrv4
    port map (
            O => \N__33435\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__6239\ : Odrv4
    port map (
            O => \N__33432\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__6238\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33424\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__33424\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\
        );

    \I__6236\ : InMux
    port map (
            O => \N__33421\,
            I => \N__33417\
        );

    \I__6235\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33414\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__33417\,
            I => \N__33411\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__33414\,
            I => \N__33408\
        );

    \I__6232\ : Odrv4
    port map (
            O => \N__33411\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__6231\ : Odrv4
    port map (
            O => \N__33408\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__6230\ : InMux
    port map (
            O => \N__33403\,
            I => \N__33400\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__33400\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\
        );

    \I__6228\ : InMux
    port map (
            O => \N__33397\,
            I => \N__33394\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__33394\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\
        );

    \I__6226\ : InMux
    port map (
            O => \N__33391\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__33388\,
            I => \N__33385\
        );

    \I__6224\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33382\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__33382\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\
        );

    \I__6222\ : InMux
    port map (
            O => \N__33379\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\
        );

    \I__6221\ : InMux
    port map (
            O => \N__33376\,
            I => \N__33373\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__33373\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\
        );

    \I__6219\ : InMux
    port map (
            O => \N__33370\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\
        );

    \I__6218\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33364\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__33364\,
            I => \N__33361\
        );

    \I__6216\ : Odrv4
    port map (
            O => \N__33361\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\
        );

    \I__6215\ : InMux
    port map (
            O => \N__33358\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\
        );

    \I__6214\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33352\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__33352\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\
        );

    \I__6212\ : InMux
    port map (
            O => \N__33349\,
            I => \bfn_14_8_0_\
        );

    \I__6211\ : InMux
    port map (
            O => \N__33346\,
            I => \N__33343\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__33343\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\
        );

    \I__6209\ : InMux
    port map (
            O => \N__33340\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\
        );

    \I__6208\ : InMux
    port map (
            O => \N__33337\,
            I => \N__33334\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__33334\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\
        );

    \I__6206\ : CascadeMux
    port map (
            O => \N__33331\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_\
        );

    \I__6205\ : InMux
    port map (
            O => \N__33328\,
            I => \N__33325\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__33325\,
            I => \N__33322\
        );

    \I__6203\ : Odrv4
    port map (
            O => \N__33322\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3\
        );

    \I__6202\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33313\
        );

    \I__6201\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33310\
        );

    \I__6200\ : InMux
    port map (
            O => \N__33317\,
            I => \N__33307\
        );

    \I__6199\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33304\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__33313\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__33310\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__33307\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__33304\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6194\ : IoInMux
    port map (
            O => \N__33295\,
            I => \N__33292\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__33292\,
            I => \N__33289\
        );

    \I__6192\ : Odrv4
    port map (
            O => \N__33289\,
            I => \current_shift_inst.timer_s1.N_180_i\
        );

    \I__6191\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33280\
        );

    \I__6190\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33280\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__33280\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\
        );

    \I__6188\ : InMux
    port map (
            O => \N__33277\,
            I => \N__33274\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__33274\,
            I => \N__33271\
        );

    \I__6186\ : Sp12to4
    port map (
            O => \N__33271\,
            I => \N__33268\
        );

    \I__6185\ : Odrv12
    port map (
            O => \N__33268\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\
        );

    \I__6184\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33262\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__33262\,
            I => \N__33259\
        );

    \I__6182\ : Span4Mux_h
    port map (
            O => \N__33259\,
            I => \N__33255\
        );

    \I__6181\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33252\
        );

    \I__6180\ : Odrv4
    port map (
            O => \N__33255\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__33252\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__6178\ : InMux
    port map (
            O => \N__33247\,
            I => \N__33244\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__33244\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\
        );

    \I__6176\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33238\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33234\
        );

    \I__6174\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33231\
        );

    \I__6173\ : Span4Mux_h
    port map (
            O => \N__33234\,
            I => \N__33228\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__33231\,
            I => \N__33225\
        );

    \I__6171\ : Odrv4
    port map (
            O => \N__33228\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__33225\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__6169\ : InMux
    port map (
            O => \N__33220\,
            I => \N__33217\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__33217\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\
        );

    \I__6167\ : InMux
    port map (
            O => \N__33214\,
            I => \N__33211\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__33211\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\
        );

    \I__6165\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33205\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__33205\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8\
        );

    \I__6163\ : CascadeMux
    port map (
            O => \N__33202\,
            I => \N__33199\
        );

    \I__6162\ : InMux
    port map (
            O => \N__33199\,
            I => \N__33195\
        );

    \I__6161\ : InMux
    port map (
            O => \N__33198\,
            I => \N__33192\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__33195\,
            I => \N__33189\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__33192\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__6158\ : Odrv4
    port map (
            O => \N__33189\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__6157\ : CascadeMux
    port map (
            O => \N__33184\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13_cascade_\
        );

    \I__6156\ : CascadeMux
    port map (
            O => \N__33181\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt19_0_cascade_\
        );

    \I__6155\ : InMux
    port map (
            O => \N__33178\,
            I => \N__33172\
        );

    \I__6154\ : InMux
    port map (
            O => \N__33177\,
            I => \N__33169\
        );

    \I__6153\ : InMux
    port map (
            O => \N__33176\,
            I => \N__33166\
        );

    \I__6152\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33163\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__33172\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__33169\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__33166\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__33163\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6147\ : CascadeMux
    port map (
            O => \N__33154\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_\
        );

    \I__6146\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33148\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__33148\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2\
        );

    \I__6144\ : InMux
    port map (
            O => \N__33145\,
            I => \N__33142\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__33142\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\
        );

    \I__6142\ : CascadeMux
    port map (
            O => \N__33139\,
            I => \N__33136\
        );

    \I__6141\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33131\
        );

    \I__6140\ : CascadeMux
    port map (
            O => \N__33135\,
            I => \N__33128\
        );

    \I__6139\ : CascadeMux
    port map (
            O => \N__33134\,
            I => \N__33125\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__33131\,
            I => \N__33122\
        );

    \I__6137\ : InMux
    port map (
            O => \N__33128\,
            I => \N__33119\
        );

    \I__6136\ : InMux
    port map (
            O => \N__33125\,
            I => \N__33116\
        );

    \I__6135\ : Span4Mux_v
    port map (
            O => \N__33122\,
            I => \N__33113\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__33119\,
            I => \N__33110\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__33116\,
            I => measured_delay_hc_19
        );

    \I__6132\ : Odrv4
    port map (
            O => \N__33113\,
            I => measured_delay_hc_19
        );

    \I__6131\ : Odrv12
    port map (
            O => \N__33110\,
            I => measured_delay_hc_19
        );

    \I__6130\ : CascadeMux
    port map (
            O => \N__33103\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__33100\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_\
        );

    \I__6128\ : CascadeMux
    port map (
            O => \N__33097\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0_cascade_\
        );

    \I__6127\ : InMux
    port map (
            O => \N__33094\,
            I => \N__33091\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__33091\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7\
        );

    \I__6125\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33085\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__33085\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0\
        );

    \I__6123\ : InMux
    port map (
            O => \N__33082\,
            I => \N__33079\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__33079\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19\
        );

    \I__6121\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33072\
        );

    \I__6120\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33069\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__33072\,
            I => \N__33062\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__33069\,
            I => \N__33062\
        );

    \I__6117\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33059\
        );

    \I__6116\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33056\
        );

    \I__6115\ : Span4Mux_v
    port map (
            O => \N__33062\,
            I => \N__33053\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__33059\,
            I => \N__33050\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__33056\,
            I => measured_delay_hc_0
        );

    \I__6112\ : Odrv4
    port map (
            O => \N__33053\,
            I => measured_delay_hc_0
        );

    \I__6111\ : Odrv4
    port map (
            O => \N__33050\,
            I => measured_delay_hc_0
        );

    \I__6110\ : InMux
    port map (
            O => \N__33043\,
            I => \N__33038\
        );

    \I__6109\ : InMux
    port map (
            O => \N__33042\,
            I => \N__33033\
        );

    \I__6108\ : InMux
    port map (
            O => \N__33041\,
            I => \N__33033\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__33038\,
            I => measured_delay_hc_20
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__33033\,
            I => measured_delay_hc_20
        );

    \I__6105\ : CascadeMux
    port map (
            O => \N__33028\,
            I => \N__33022\
        );

    \I__6104\ : InMux
    port map (
            O => \N__33027\,
            I => \N__33018\
        );

    \I__6103\ : InMux
    port map (
            O => \N__33026\,
            I => \N__33015\
        );

    \I__6102\ : InMux
    port map (
            O => \N__33025\,
            I => \N__33010\
        );

    \I__6101\ : InMux
    port map (
            O => \N__33022\,
            I => \N__33010\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__33021\,
            I => \N__33007\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__33018\,
            I => \N__33004\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__33015\,
            I => \N__32999\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__33010\,
            I => \N__32999\
        );

    \I__6096\ : InMux
    port map (
            O => \N__33007\,
            I => \N__32996\
        );

    \I__6095\ : Span4Mux_h
    port map (
            O => \N__33004\,
            I => \N__32993\
        );

    \I__6094\ : Span4Mux_h
    port map (
            O => \N__32999\,
            I => \N__32990\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__32996\,
            I => measured_delay_hc_16
        );

    \I__6092\ : Odrv4
    port map (
            O => \N__32993\,
            I => measured_delay_hc_16
        );

    \I__6091\ : Odrv4
    port map (
            O => \N__32990\,
            I => measured_delay_hc_16
        );

    \I__6090\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32978\
        );

    \I__6089\ : InMux
    port map (
            O => \N__32982\,
            I => \N__32975\
        );

    \I__6088\ : CascadeMux
    port map (
            O => \N__32981\,
            I => \N__32971\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__32978\,
            I => \N__32966\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32966\
        );

    \I__6085\ : InMux
    port map (
            O => \N__32974\,
            I => \N__32963\
        );

    \I__6084\ : InMux
    port map (
            O => \N__32971\,
            I => \N__32960\
        );

    \I__6083\ : Span4Mux_h
    port map (
            O => \N__32966\,
            I => \N__32957\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__32963\,
            I => \N__32954\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__32960\,
            I => measured_delay_hc_1
        );

    \I__6080\ : Odrv4
    port map (
            O => \N__32957\,
            I => measured_delay_hc_1
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__32954\,
            I => measured_delay_hc_1
        );

    \I__6078\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32943\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32940\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__32943\,
            I => \N__32935\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__32940\,
            I => \N__32932\
        );

    \I__6074\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32929\
        );

    \I__6073\ : InMux
    port map (
            O => \N__32938\,
            I => \N__32926\
        );

    \I__6072\ : Span4Mux_h
    port map (
            O => \N__32935\,
            I => \N__32923\
        );

    \I__6071\ : Span4Mux_v
    port map (
            O => \N__32932\,
            I => \N__32918\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__32929\,
            I => \N__32918\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__32926\,
            I => measured_delay_hc_8
        );

    \I__6068\ : Odrv4
    port map (
            O => \N__32923\,
            I => measured_delay_hc_8
        );

    \I__6067\ : Odrv4
    port map (
            O => \N__32918\,
            I => measured_delay_hc_8
        );

    \I__6066\ : InMux
    port map (
            O => \N__32911\,
            I => \N__32904\
        );

    \I__6065\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32904\
        );

    \I__6064\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32901\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__32904\,
            I => \N__32898\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__32901\,
            I => measured_delay_hc_21
        );

    \I__6061\ : Odrv4
    port map (
            O => \N__32898\,
            I => measured_delay_hc_21
        );

    \I__6060\ : InMux
    port map (
            O => \N__32893\,
            I => \N__32886\
        );

    \I__6059\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32883\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32880\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32890\,
            I => \N__32877\
        );

    \I__6056\ : CascadeMux
    port map (
            O => \N__32889\,
            I => \N__32874\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__32886\,
            I => \N__32871\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__32883\,
            I => \N__32868\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__32880\,
            I => \N__32865\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__32877\,
            I => \N__32862\
        );

    \I__6051\ : InMux
    port map (
            O => \N__32874\,
            I => \N__32859\
        );

    \I__6050\ : Span4Mux_h
    port map (
            O => \N__32871\,
            I => \N__32856\
        );

    \I__6049\ : Span4Mux_v
    port map (
            O => \N__32868\,
            I => \N__32851\
        );

    \I__6048\ : Span4Mux_v
    port map (
            O => \N__32865\,
            I => \N__32851\
        );

    \I__6047\ : Span4Mux_h
    port map (
            O => \N__32862\,
            I => \N__32848\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__32859\,
            I => measured_delay_hc_15
        );

    \I__6045\ : Odrv4
    port map (
            O => \N__32856\,
            I => measured_delay_hc_15
        );

    \I__6044\ : Odrv4
    port map (
            O => \N__32851\,
            I => measured_delay_hc_15
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__32848\,
            I => measured_delay_hc_15
        );

    \I__6042\ : InMux
    port map (
            O => \N__32839\,
            I => \N__32836\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__32836\,
            I => \N__32831\
        );

    \I__6040\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32828\
        );

    \I__6039\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32824\
        );

    \I__6038\ : Span4Mux_h
    port map (
            O => \N__32831\,
            I => \N__32818\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__32828\,
            I => \N__32818\
        );

    \I__6036\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32815\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__32824\,
            I => \N__32812\
        );

    \I__6034\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32809\
        );

    \I__6033\ : Span4Mux_v
    port map (
            O => \N__32818\,
            I => \N__32802\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__32815\,
            I => \N__32802\
        );

    \I__6031\ : Span4Mux_h
    port map (
            O => \N__32812\,
            I => \N__32802\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__32809\,
            I => measured_delay_hc_4
        );

    \I__6029\ : Odrv4
    port map (
            O => \N__32802\,
            I => measured_delay_hc_4
        );

    \I__6028\ : CascadeMux
    port map (
            O => \N__32797\,
            I => \N__32793\
        );

    \I__6027\ : CascadeMux
    port map (
            O => \N__32796\,
            I => \N__32790\
        );

    \I__6026\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32787\
        );

    \I__6025\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32784\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__32787\,
            I => \N__32779\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__32784\,
            I => \N__32779\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__32779\,
            I => \N__32774\
        );

    \I__6021\ : InMux
    port map (
            O => \N__32778\,
            I => \N__32771\
        );

    \I__6020\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32768\
        );

    \I__6019\ : Sp12to4
    port map (
            O => \N__32774\,
            I => \N__32763\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__32771\,
            I => \N__32763\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__32768\,
            I => measured_delay_hc_2
        );

    \I__6016\ : Odrv12
    port map (
            O => \N__32763\,
            I => measured_delay_hc_2
        );

    \I__6015\ : InMux
    port map (
            O => \N__32758\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__6014\ : InMux
    port map (
            O => \N__32755\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__6013\ : InMux
    port map (
            O => \N__32752\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32749\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__6011\ : InMux
    port map (
            O => \N__32746\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__6010\ : InMux
    port map (
            O => \N__32743\,
            I => \N__32737\
        );

    \I__6009\ : InMux
    port map (
            O => \N__32742\,
            I => \N__32737\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__32737\,
            I => \N__32734\
        );

    \I__6007\ : Odrv4
    port map (
            O => \N__32734\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt3\
        );

    \I__6006\ : InMux
    port map (
            O => \N__32731\,
            I => \N__32727\
        );

    \I__6005\ : InMux
    port map (
            O => \N__32730\,
            I => \N__32724\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__32727\,
            I => \N__32721\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__32724\,
            I => \N__32718\
        );

    \I__6002\ : Span4Mux_h
    port map (
            O => \N__32721\,
            I => \N__32714\
        );

    \I__6001\ : Span4Mux_h
    port map (
            O => \N__32718\,
            I => \N__32711\
        );

    \I__6000\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32708\
        );

    \I__5999\ : Odrv4
    port map (
            O => \N__32714\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__5998\ : Odrv4
    port map (
            O => \N__32711\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__32708\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__5996\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32698\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__32698\,
            I => \N__32695\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__32695\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__32692\,
            I => \N__32687\
        );

    \I__5992\ : InMux
    port map (
            O => \N__32691\,
            I => \N__32684\
        );

    \I__5991\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32679\
        );

    \I__5990\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32679\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__32684\,
            I => measured_delay_hc_22
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__32679\,
            I => measured_delay_hc_22
        );

    \I__5987\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32669\
        );

    \I__5986\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32666\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__32672\,
            I => \N__32663\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__32669\,
            I => \N__32660\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__32666\,
            I => \N__32657\
        );

    \I__5982\ : InMux
    port map (
            O => \N__32663\,
            I => \N__32653\
        );

    \I__5981\ : Span4Mux_v
    port map (
            O => \N__32660\,
            I => \N__32650\
        );

    \I__5980\ : Span4Mux_h
    port map (
            O => \N__32657\,
            I => \N__32647\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32644\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__32653\,
            I => measured_delay_hc_7
        );

    \I__5977\ : Odrv4
    port map (
            O => \N__32650\,
            I => measured_delay_hc_7
        );

    \I__5976\ : Odrv4
    port map (
            O => \N__32647\,
            I => measured_delay_hc_7
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__32644\,
            I => measured_delay_hc_7
        );

    \I__5974\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32632\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__32632\,
            I => \N__32629\
        );

    \I__5972\ : Span4Mux_v
    port map (
            O => \N__32629\,
            I => \N__32626\
        );

    \I__5971\ : Odrv4
    port map (
            O => \N__32626\,
            I => \current_shift_inst.un38_control_input_0_s0_19\
        );

    \I__5970\ : InMux
    port map (
            O => \N__32623\,
            I => \current_shift_inst.un38_control_input_cry_18_s0\
        );

    \I__5969\ : InMux
    port map (
            O => \N__32620\,
            I => \N__32617\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__32617\,
            I => \N__32614\
        );

    \I__5967\ : Odrv12
    port map (
            O => \N__32614\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__5966\ : InMux
    port map (
            O => \N__32611\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__5965\ : InMux
    port map (
            O => \N__32608\,
            I => \N__32605\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__32605\,
            I => \N__32602\
        );

    \I__5963\ : Odrv12
    port map (
            O => \N__32602\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__5962\ : InMux
    port map (
            O => \N__32599\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__5961\ : CascadeMux
    port map (
            O => \N__32596\,
            I => \N__32593\
        );

    \I__5960\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32590\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__32590\,
            I => \N__32587\
        );

    \I__5958\ : Odrv12
    port map (
            O => \N__32587\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__5957\ : InMux
    port map (
            O => \N__32584\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__5956\ : InMux
    port map (
            O => \N__32581\,
            I => \N__32578\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__32578\,
            I => \N__32575\
        );

    \I__5954\ : Odrv12
    port map (
            O => \N__32575\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__5953\ : InMux
    port map (
            O => \N__32572\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__5952\ : InMux
    port map (
            O => \N__32569\,
            I => \bfn_13_20_0_\
        );

    \I__5951\ : InMux
    port map (
            O => \N__32566\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__5950\ : InMux
    port map (
            O => \N__32563\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__5949\ : InMux
    port map (
            O => \N__32560\,
            I => \current_shift_inst.un38_control_input_cry_9_s0\
        );

    \I__5948\ : InMux
    port map (
            O => \N__32557\,
            I => \current_shift_inst.un38_control_input_cry_10_s0\
        );

    \I__5947\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32551\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__32551\,
            I => \N__32548\
        );

    \I__5945\ : Odrv12
    port map (
            O => \N__32548\,
            I => \current_shift_inst.un38_control_input_0_s0_12\
        );

    \I__5944\ : InMux
    port map (
            O => \N__32545\,
            I => \current_shift_inst.un38_control_input_cry_11_s0\
        );

    \I__5943\ : InMux
    port map (
            O => \N__32542\,
            I => \N__32539\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__32539\,
            I => \N__32536\
        );

    \I__5941\ : Odrv12
    port map (
            O => \N__32536\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\
        );

    \I__5940\ : InMux
    port map (
            O => \N__32533\,
            I => \current_shift_inst.un38_control_input_cry_12_s0\
        );

    \I__5939\ : InMux
    port map (
            O => \N__32530\,
            I => \N__32527\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__32527\,
            I => \N__32524\
        );

    \I__5937\ : Odrv4
    port map (
            O => \N__32524\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\
        );

    \I__5936\ : InMux
    port map (
            O => \N__32521\,
            I => \N__32518\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__32518\,
            I => \N__32515\
        );

    \I__5934\ : Odrv12
    port map (
            O => \N__32515\,
            I => \current_shift_inst.un38_control_input_0_s0_14\
        );

    \I__5933\ : InMux
    port map (
            O => \N__32512\,
            I => \current_shift_inst.un38_control_input_cry_13_s0\
        );

    \I__5932\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32506\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__32506\,
            I => \N__32503\
        );

    \I__5930\ : Odrv12
    port map (
            O => \N__32503\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\
        );

    \I__5929\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32497\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__32497\,
            I => \N__32494\
        );

    \I__5927\ : Odrv4
    port map (
            O => \N__32494\,
            I => \current_shift_inst.un38_control_input_0_s0_15\
        );

    \I__5926\ : InMux
    port map (
            O => \N__32491\,
            I => \current_shift_inst.un38_control_input_cry_14_s0\
        );

    \I__5925\ : InMux
    port map (
            O => \N__32488\,
            I => \N__32485\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__32485\,
            I => \N__32482\
        );

    \I__5923\ : Span4Mux_v
    port map (
            O => \N__32482\,
            I => \N__32479\
        );

    \I__5922\ : Odrv4
    port map (
            O => \N__32479\,
            I => \current_shift_inst.un38_control_input_0_s0_16\
        );

    \I__5921\ : InMux
    port map (
            O => \N__32476\,
            I => \bfn_13_19_0_\
        );

    \I__5920\ : InMux
    port map (
            O => \N__32473\,
            I => \N__32470\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__32470\,
            I => \N__32467\
        );

    \I__5918\ : Span4Mux_h
    port map (
            O => \N__32467\,
            I => \N__32464\
        );

    \I__5917\ : Odrv4
    port map (
            O => \N__32464\,
            I => \current_shift_inst.un38_control_input_0_s0_17\
        );

    \I__5916\ : InMux
    port map (
            O => \N__32461\,
            I => \current_shift_inst.un38_control_input_cry_16_s0\
        );

    \I__5915\ : InMux
    port map (
            O => \N__32458\,
            I => \N__32455\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__32455\,
            I => \N__32452\
        );

    \I__5913\ : Odrv12
    port map (
            O => \N__32452\,
            I => \current_shift_inst.un38_control_input_0_s0_18\
        );

    \I__5912\ : InMux
    port map (
            O => \N__32449\,
            I => \current_shift_inst.un38_control_input_cry_17_s0\
        );

    \I__5911\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32443\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__32443\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__5909\ : InMux
    port map (
            O => \N__32440\,
            I => \N__32437\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__32437\,
            I => \N__32434\
        );

    \I__5907\ : Odrv4
    port map (
            O => \N__32434\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__5906\ : InMux
    port map (
            O => \N__32431\,
            I => \current_shift_inst.un38_control_input_cry_5_s0\
        );

    \I__5905\ : InMux
    port map (
            O => \N__32428\,
            I => \N__32425\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__32425\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\
        );

    \I__5903\ : InMux
    port map (
            O => \N__32422\,
            I => \current_shift_inst.un38_control_input_cry_6_s0\
        );

    \I__5902\ : InMux
    port map (
            O => \N__32419\,
            I => \N__32416\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__32416\,
            I => \N__32413\
        );

    \I__5900\ : Odrv4
    port map (
            O => \N__32413\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\
        );

    \I__5899\ : InMux
    port map (
            O => \N__32410\,
            I => \N__32407\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__32407\,
            I => \N__32404\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__32404\,
            I => \current_shift_inst.un38_control_input_0_s0_8\
        );

    \I__5896\ : InMux
    port map (
            O => \N__32401\,
            I => \bfn_13_18_0_\
        );

    \I__5895\ : InMux
    port map (
            O => \N__32398\,
            I => \N__32395\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__32395\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\
        );

    \I__5893\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32389\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__32389\,
            I => \N__32386\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__32386\,
            I => \current_shift_inst.un38_control_input_0_s0_9\
        );

    \I__5890\ : InMux
    port map (
            O => \N__32383\,
            I => \current_shift_inst.un38_control_input_cry_8_s0\
        );

    \I__5889\ : InMux
    port map (
            O => \N__32380\,
            I => \N__32377\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__32377\,
            I => \N__32374\
        );

    \I__5887\ : Odrv4
    port map (
            O => \N__32374\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\
        );

    \I__5886\ : InMux
    port map (
            O => \N__32371\,
            I => \N__32368\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__32368\,
            I => \N__32365\
        );

    \I__5884\ : Odrv4
    port map (
            O => \N__32365\,
            I => \current_shift_inst.un38_control_input_0_s0_10\
        );

    \I__5883\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32359\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__32359\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__5881\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32353\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__32353\,
            I => \N__32350\
        );

    \I__5879\ : Odrv12
    port map (
            O => \N__32350\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__5878\ : InMux
    port map (
            O => \N__32347\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_24\
        );

    \I__5877\ : InMux
    port map (
            O => \N__32344\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_25\
        );

    \I__5876\ : InMux
    port map (
            O => \N__32341\,
            I => \N__32338\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__32338\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\
        );

    \I__5874\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32332\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__32332\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\
        );

    \I__5872\ : InMux
    port map (
            O => \N__32329\,
            I => \N__32326\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__32326\,
            I => \N__32323\
        );

    \I__5870\ : Odrv4
    port map (
            O => \N__32323\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\
        );

    \I__5869\ : InMux
    port map (
            O => \N__32320\,
            I => \bfn_13_12_0_\
        );

    \I__5868\ : InMux
    port map (
            O => \N__32317\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_16\
        );

    \I__5867\ : InMux
    port map (
            O => \N__32314\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_17\
        );

    \I__5866\ : InMux
    port map (
            O => \N__32311\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_18\
        );

    \I__5865\ : InMux
    port map (
            O => \N__32308\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_19\
        );

    \I__5864\ : InMux
    port map (
            O => \N__32305\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_20\
        );

    \I__5863\ : InMux
    port map (
            O => \N__32302\,
            I => \N__32299\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__32299\,
            I => \N__32296\
        );

    \I__5861\ : Span4Mux_v
    port map (
            O => \N__32296\,
            I => \N__32293\
        );

    \I__5860\ : Odrv4
    port map (
            O => \N__32293\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\
        );

    \I__5859\ : InMux
    port map (
            O => \N__32290\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_21\
        );

    \I__5858\ : InMux
    port map (
            O => \N__32287\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_22\
        );

    \I__5857\ : InMux
    port map (
            O => \N__32284\,
            I => \bfn_13_13_0_\
        );

    \I__5856\ : InMux
    port map (
            O => \N__32281\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__5855\ : InMux
    port map (
            O => \N__32278\,
            I => \bfn_13_11_0_\
        );

    \I__5854\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32272\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__32272\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__5852\ : InMux
    port map (
            O => \N__32269\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__5851\ : InMux
    port map (
            O => \N__32266\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__5850\ : InMux
    port map (
            O => \N__32263\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__5849\ : InMux
    port map (
            O => \N__32260\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__5848\ : InMux
    port map (
            O => \N__32257\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__5847\ : InMux
    port map (
            O => \N__32254\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__5846\ : InMux
    port map (
            O => \N__32251\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_14\
        );

    \I__5845\ : InMux
    port map (
            O => \N__32248\,
            I => \N__32245\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__32245\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__5843\ : InMux
    port map (
            O => \N__32242\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__5842\ : InMux
    port map (
            O => \N__32239\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__5841\ : InMux
    port map (
            O => \N__32236\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__5840\ : InMux
    port map (
            O => \N__32233\,
            I => \N__32230\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__32230\,
            I => \N__32227\
        );

    \I__5838\ : Span4Mux_h
    port map (
            O => \N__32227\,
            I => \N__32224\
        );

    \I__5837\ : Odrv4
    port map (
            O => \N__32224\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__5836\ : InMux
    port map (
            O => \N__32221\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__5835\ : InMux
    port map (
            O => \N__32218\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__5834\ : InMux
    port map (
            O => \N__32215\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__32212\,
            I => \N__32208\
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__32211\,
            I => \N__32205\
        );

    \I__5831\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32202\
        );

    \I__5830\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32198\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__32202\,
            I => \N__32195\
        );

    \I__5828\ : InMux
    port map (
            O => \N__32201\,
            I => \N__32192\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__32198\,
            I => \N__32188\
        );

    \I__5826\ : Span4Mux_h
    port map (
            O => \N__32195\,
            I => \N__32183\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__32192\,
            I => \N__32183\
        );

    \I__5824\ : InMux
    port map (
            O => \N__32191\,
            I => \N__32180\
        );

    \I__5823\ : Span4Mux_h
    port map (
            O => \N__32188\,
            I => \N__32177\
        );

    \I__5822\ : Span4Mux_v
    port map (
            O => \N__32183\,
            I => \N__32174\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__32180\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5820\ : Odrv4
    port map (
            O => \N__32177\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5819\ : Odrv4
    port map (
            O => \N__32174\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5818\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32163\
        );

    \I__5817\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32160\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__32163\,
            I => measured_delay_hc_23
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__32160\,
            I => measured_delay_hc_23
        );

    \I__5814\ : InMux
    port map (
            O => \N__32155\,
            I => \N__32151\
        );

    \I__5813\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32148\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__32151\,
            I => \N__32144\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__32148\,
            I => \N__32141\
        );

    \I__5810\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32138\
        );

    \I__5809\ : Span4Mux_s3_v
    port map (
            O => \N__32144\,
            I => \N__32135\
        );

    \I__5808\ : Span4Mux_s3_v
    port map (
            O => \N__32141\,
            I => \N__32132\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__32138\,
            I => \N__32129\
        );

    \I__5806\ : Span4Mux_v
    port map (
            O => \N__32135\,
            I => \N__32126\
        );

    \I__5805\ : Span4Mux_v
    port map (
            O => \N__32132\,
            I => \N__32123\
        );

    \I__5804\ : Span12Mux_h
    port map (
            O => \N__32129\,
            I => \N__32117\
        );

    \I__5803\ : Sp12to4
    port map (
            O => \N__32126\,
            I => \N__32112\
        );

    \I__5802\ : Sp12to4
    port map (
            O => \N__32123\,
            I => \N__32112\
        );

    \I__5801\ : InMux
    port map (
            O => \N__32122\,
            I => \N__32109\
        );

    \I__5800\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32104\
        );

    \I__5799\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32104\
        );

    \I__5798\ : Span12Mux_v
    port map (
            O => \N__32117\,
            I => \N__32101\
        );

    \I__5797\ : Span12Mux_h
    port map (
            O => \N__32112\,
            I => \N__32096\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__32109\,
            I => \N__32096\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__32104\,
            I => state_3
        );

    \I__5794\ : Odrv12
    port map (
            O => \N__32101\,
            I => state_3
        );

    \I__5793\ : Odrv12
    port map (
            O => \N__32096\,
            I => state_3
        );

    \I__5792\ : IoInMux
    port map (
            O => \N__32089\,
            I => \N__32086\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__32086\,
            I => \N__32083\
        );

    \I__5790\ : Span4Mux_s2_v
    port map (
            O => \N__32083\,
            I => \N__32079\
        );

    \I__5789\ : CascadeMux
    port map (
            O => \N__32082\,
            I => \N__32076\
        );

    \I__5788\ : Span4Mux_h
    port map (
            O => \N__32079\,
            I => \N__32072\
        );

    \I__5787\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32069\
        );

    \I__5786\ : InMux
    port map (
            O => \N__32075\,
            I => \N__32066\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__32072\,
            I => s1_phy_c
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__32069\,
            I => s1_phy_c
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__32066\,
            I => s1_phy_c
        );

    \I__5782\ : CascadeMux
    port map (
            O => \N__32059\,
            I => \N__32056\
        );

    \I__5781\ : InMux
    port map (
            O => \N__32056\,
            I => \N__32053\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__32053\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__32050\,
            I => \current_shift_inst.PI_CTRL.un1_enablelt3_0_cascade_\
        );

    \I__5778\ : InMux
    port map (
            O => \N__32047\,
            I => \N__32044\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__32044\,
            I => \N__32041\
        );

    \I__5776\ : Odrv4
    port map (
            O => \N__32041\,
            I => \current_shift_inst.PI_CTRL.N_71\
        );

    \I__5775\ : CascadeMux
    port map (
            O => \N__32038\,
            I => \N__32031\
        );

    \I__5774\ : InMux
    port map (
            O => \N__32037\,
            I => \N__32028\
        );

    \I__5773\ : InMux
    port map (
            O => \N__32036\,
            I => \N__32025\
        );

    \I__5772\ : InMux
    port map (
            O => \N__32035\,
            I => \N__32020\
        );

    \I__5771\ : InMux
    port map (
            O => \N__32034\,
            I => \N__32020\
        );

    \I__5770\ : InMux
    port map (
            O => \N__32031\,
            I => \N__32017\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__32028\,
            I => \N__32014\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__32025\,
            I => \N__32009\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__32020\,
            I => \N__32009\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__32017\,
            I => measured_delay_hc_11
        );

    \I__5765\ : Odrv12
    port map (
            O => \N__32014\,
            I => measured_delay_hc_11
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__32009\,
            I => measured_delay_hc_11
        );

    \I__5763\ : CascadeMux
    port map (
            O => \N__32002\,
            I => \N__31997\
        );

    \I__5762\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31993\
        );

    \I__5761\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31987\
        );

    \I__5760\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31987\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__31996\,
            I => \N__31984\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__31993\,
            I => \N__31981\
        );

    \I__5757\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31978\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__31987\,
            I => \N__31975\
        );

    \I__5755\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31972\
        );

    \I__5754\ : Span12Mux_v
    port map (
            O => \N__31981\,
            I => \N__31969\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__31978\,
            I => \N__31964\
        );

    \I__5752\ : Span4Mux_h
    port map (
            O => \N__31975\,
            I => \N__31964\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__31972\,
            I => measured_delay_hc_9
        );

    \I__5750\ : Odrv12
    port map (
            O => \N__31969\,
            I => measured_delay_hc_9
        );

    \I__5749\ : Odrv4
    port map (
            O => \N__31964\,
            I => measured_delay_hc_9
        );

    \I__5748\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31954\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__31954\,
            I => \N__31948\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__31953\,
            I => \N__31945\
        );

    \I__5745\ : InMux
    port map (
            O => \N__31952\,
            I => \N__31942\
        );

    \I__5744\ : CascadeMux
    port map (
            O => \N__31951\,
            I => \N__31938\
        );

    \I__5743\ : Span4Mux_h
    port map (
            O => \N__31948\,
            I => \N__31935\
        );

    \I__5742\ : InMux
    port map (
            O => \N__31945\,
            I => \N__31932\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__31942\,
            I => \N__31929\
        );

    \I__5740\ : InMux
    port map (
            O => \N__31941\,
            I => \N__31926\
        );

    \I__5739\ : InMux
    port map (
            O => \N__31938\,
            I => \N__31923\
        );

    \I__5738\ : Span4Mux_v
    port map (
            O => \N__31935\,
            I => \N__31920\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__31932\,
            I => \N__31915\
        );

    \I__5736\ : Span4Mux_h
    port map (
            O => \N__31929\,
            I => \N__31915\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__31926\,
            I => \N__31912\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__31923\,
            I => measured_delay_hc_14
        );

    \I__5733\ : Odrv4
    port map (
            O => \N__31920\,
            I => measured_delay_hc_14
        );

    \I__5732\ : Odrv4
    port map (
            O => \N__31915\,
            I => measured_delay_hc_14
        );

    \I__5731\ : Odrv12
    port map (
            O => \N__31912\,
            I => measured_delay_hc_14
        );

    \I__5730\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31898\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__31902\,
            I => \N__31894\
        );

    \I__5728\ : CascadeMux
    port map (
            O => \N__31901\,
            I => \N__31891\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__31898\,
            I => \N__31888\
        );

    \I__5726\ : InMux
    port map (
            O => \N__31897\,
            I => \N__31885\
        );

    \I__5725\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31880\
        );

    \I__5724\ : InMux
    port map (
            O => \N__31891\,
            I => \N__31880\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__31888\,
            I => \N__31876\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__31885\,
            I => \N__31873\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__31880\,
            I => \N__31870\
        );

    \I__5720\ : InMux
    port map (
            O => \N__31879\,
            I => \N__31867\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__31876\,
            I => \N__31864\
        );

    \I__5718\ : Span4Mux_h
    port map (
            O => \N__31873\,
            I => \N__31859\
        );

    \I__5717\ : Span4Mux_h
    port map (
            O => \N__31870\,
            I => \N__31859\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__31867\,
            I => measured_delay_hc_6
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__31864\,
            I => measured_delay_hc_6
        );

    \I__5714\ : Odrv4
    port map (
            O => \N__31859\,
            I => measured_delay_hc_6
        );

    \I__5713\ : InMux
    port map (
            O => \N__31852\,
            I => \N__31845\
        );

    \I__5712\ : InMux
    port map (
            O => \N__31851\,
            I => \N__31842\
        );

    \I__5711\ : InMux
    port map (
            O => \N__31850\,
            I => \N__31839\
        );

    \I__5710\ : CascadeMux
    port map (
            O => \N__31849\,
            I => \N__31836\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__31848\,
            I => \N__31833\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__31845\,
            I => \N__31830\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__31842\,
            I => \N__31825\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__31839\,
            I => \N__31825\
        );

    \I__5705\ : InMux
    port map (
            O => \N__31836\,
            I => \N__31822\
        );

    \I__5704\ : InMux
    port map (
            O => \N__31833\,
            I => \N__31819\
        );

    \I__5703\ : Span12Mux_h
    port map (
            O => \N__31830\,
            I => \N__31812\
        );

    \I__5702\ : Sp12to4
    port map (
            O => \N__31825\,
            I => \N__31812\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__31822\,
            I => \N__31812\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__31819\,
            I => measured_delay_hc_13
        );

    \I__5699\ : Odrv12
    port map (
            O => \N__31812\,
            I => measured_delay_hc_13
        );

    \I__5698\ : InMux
    port map (
            O => \N__31807\,
            I => \N__31803\
        );

    \I__5697\ : InMux
    port map (
            O => \N__31806\,
            I => \N__31800\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__31803\,
            I => measured_delay_hc_24
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__31800\,
            I => measured_delay_hc_24
        );

    \I__5694\ : InMux
    port map (
            O => \N__31795\,
            I => \N__31791\
        );

    \I__5693\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31788\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__31791\,
            I => measured_delay_hc_25
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__31788\,
            I => measured_delay_hc_25
        );

    \I__5690\ : CascadeMux
    port map (
            O => \N__31783\,
            I => \N__31779\
        );

    \I__5689\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31776\
        );

    \I__5688\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31773\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__31776\,
            I => measured_delay_hc_26
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__31773\,
            I => measured_delay_hc_26
        );

    \I__5685\ : CascadeMux
    port map (
            O => \N__31768\,
            I => \N__31765\
        );

    \I__5684\ : InMux
    port map (
            O => \N__31765\,
            I => \N__31762\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__31762\,
            I => \N__31759\
        );

    \I__5682\ : Odrv4
    port map (
            O => \N__31759\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__5681\ : InMux
    port map (
            O => \N__31756\,
            I => \N__31720\
        );

    \I__5680\ : InMux
    port map (
            O => \N__31755\,
            I => \N__31720\
        );

    \I__5679\ : InMux
    port map (
            O => \N__31754\,
            I => \N__31720\
        );

    \I__5678\ : InMux
    port map (
            O => \N__31753\,
            I => \N__31720\
        );

    \I__5677\ : InMux
    port map (
            O => \N__31752\,
            I => \N__31720\
        );

    \I__5676\ : InMux
    port map (
            O => \N__31751\,
            I => \N__31704\
        );

    \I__5675\ : InMux
    port map (
            O => \N__31750\,
            I => \N__31704\
        );

    \I__5674\ : InMux
    port map (
            O => \N__31749\,
            I => \N__31704\
        );

    \I__5673\ : InMux
    port map (
            O => \N__31748\,
            I => \N__31704\
        );

    \I__5672\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31704\
        );

    \I__5671\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31689\
        );

    \I__5670\ : InMux
    port map (
            O => \N__31745\,
            I => \N__31689\
        );

    \I__5669\ : InMux
    port map (
            O => \N__31744\,
            I => \N__31689\
        );

    \I__5668\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31689\
        );

    \I__5667\ : InMux
    port map (
            O => \N__31742\,
            I => \N__31689\
        );

    \I__5666\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31689\
        );

    \I__5665\ : InMux
    port map (
            O => \N__31740\,
            I => \N__31689\
        );

    \I__5664\ : InMux
    port map (
            O => \N__31739\,
            I => \N__31678\
        );

    \I__5663\ : InMux
    port map (
            O => \N__31738\,
            I => \N__31678\
        );

    \I__5662\ : InMux
    port map (
            O => \N__31737\,
            I => \N__31678\
        );

    \I__5661\ : InMux
    port map (
            O => \N__31736\,
            I => \N__31678\
        );

    \I__5660\ : InMux
    port map (
            O => \N__31735\,
            I => \N__31678\
        );

    \I__5659\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31669\
        );

    \I__5658\ : InMux
    port map (
            O => \N__31733\,
            I => \N__31669\
        );

    \I__5657\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31669\
        );

    \I__5656\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31669\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__31720\,
            I => \N__31659\
        );

    \I__5654\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31648\
        );

    \I__5653\ : InMux
    port map (
            O => \N__31718\,
            I => \N__31648\
        );

    \I__5652\ : InMux
    port map (
            O => \N__31717\,
            I => \N__31648\
        );

    \I__5651\ : InMux
    port map (
            O => \N__31716\,
            I => \N__31648\
        );

    \I__5650\ : InMux
    port map (
            O => \N__31715\,
            I => \N__31648\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__31704\,
            I => \N__31643\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__31689\,
            I => \N__31643\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__31678\,
            I => \N__31638\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__31669\,
            I => \N__31638\
        );

    \I__5645\ : InMux
    port map (
            O => \N__31668\,
            I => \N__31629\
        );

    \I__5644\ : InMux
    port map (
            O => \N__31667\,
            I => \N__31629\
        );

    \I__5643\ : InMux
    port map (
            O => \N__31666\,
            I => \N__31629\
        );

    \I__5642\ : InMux
    port map (
            O => \N__31665\,
            I => \N__31629\
        );

    \I__5641\ : InMux
    port map (
            O => \N__31664\,
            I => \N__31622\
        );

    \I__5640\ : InMux
    port map (
            O => \N__31663\,
            I => \N__31622\
        );

    \I__5639\ : InMux
    port map (
            O => \N__31662\,
            I => \N__31622\
        );

    \I__5638\ : Odrv4
    port map (
            O => \N__31659\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__31648\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__5636\ : Odrv4
    port map (
            O => \N__31643\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__5635\ : Odrv4
    port map (
            O => \N__31638\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__31629\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__31622\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__31609\,
            I => \N__31606\
        );

    \I__5631\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31603\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__31603\,
            I => \N__31600\
        );

    \I__5629\ : Span4Mux_h
    port map (
            O => \N__31600\,
            I => \N__31597\
        );

    \I__5628\ : Odrv4
    port map (
            O => \N__31597\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__5627\ : CEMux
    port map (
            O => \N__31594\,
            I => \N__31591\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__31591\,
            I => \N__31588\
        );

    \I__5625\ : Span4Mux_h
    port map (
            O => \N__31588\,
            I => \N__31585\
        );

    \I__5624\ : Span4Mux_h
    port map (
            O => \N__31585\,
            I => \N__31579\
        );

    \I__5623\ : CEMux
    port map (
            O => \N__31584\,
            I => \N__31576\
        );

    \I__5622\ : CEMux
    port map (
            O => \N__31583\,
            I => \N__31573\
        );

    \I__5621\ : CEMux
    port map (
            O => \N__31582\,
            I => \N__31570\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__31579\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__31576\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__31573\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__31570\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5616\ : CascadeMux
    port map (
            O => \N__31561\,
            I => \N__31555\
        );

    \I__5615\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31552\
        );

    \I__5614\ : InMux
    port map (
            O => \N__31559\,
            I => \N__31546\
        );

    \I__5613\ : InMux
    port map (
            O => \N__31558\,
            I => \N__31546\
        );

    \I__5612\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31543\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__31552\,
            I => \N__31540\
        );

    \I__5610\ : InMux
    port map (
            O => \N__31551\,
            I => \N__31537\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__31546\,
            I => \N__31534\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__31543\,
            I => measured_delay_hc_10
        );

    \I__5607\ : Odrv12
    port map (
            O => \N__31540\,
            I => measured_delay_hc_10
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__31537\,
            I => measured_delay_hc_10
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__31534\,
            I => measured_delay_hc_10
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__31525\,
            I => \N__31517\
        );

    \I__5603\ : CascadeMux
    port map (
            O => \N__31524\,
            I => \N__31514\
        );

    \I__5602\ : CascadeMux
    port map (
            O => \N__31523\,
            I => \N__31503\
        );

    \I__5601\ : CascadeMux
    port map (
            O => \N__31522\,
            I => \N__31494\
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__31521\,
            I => \N__31489\
        );

    \I__5599\ : CascadeMux
    port map (
            O => \N__31520\,
            I => \N__31486\
        );

    \I__5598\ : InMux
    port map (
            O => \N__31517\,
            I => \N__31467\
        );

    \I__5597\ : InMux
    port map (
            O => \N__31514\,
            I => \N__31467\
        );

    \I__5596\ : InMux
    port map (
            O => \N__31513\,
            I => \N__31467\
        );

    \I__5595\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31467\
        );

    \I__5594\ : InMux
    port map (
            O => \N__31511\,
            I => \N__31467\
        );

    \I__5593\ : InMux
    port map (
            O => \N__31510\,
            I => \N__31456\
        );

    \I__5592\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31456\
        );

    \I__5591\ : InMux
    port map (
            O => \N__31508\,
            I => \N__31456\
        );

    \I__5590\ : InMux
    port map (
            O => \N__31507\,
            I => \N__31456\
        );

    \I__5589\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31456\
        );

    \I__5588\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31441\
        );

    \I__5587\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31441\
        );

    \I__5586\ : InMux
    port map (
            O => \N__31501\,
            I => \N__31441\
        );

    \I__5585\ : InMux
    port map (
            O => \N__31500\,
            I => \N__31441\
        );

    \I__5584\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31441\
        );

    \I__5583\ : InMux
    port map (
            O => \N__31498\,
            I => \N__31441\
        );

    \I__5582\ : InMux
    port map (
            O => \N__31497\,
            I => \N__31441\
        );

    \I__5581\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31437\
        );

    \I__5580\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31428\
        );

    \I__5579\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31428\
        );

    \I__5578\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31428\
        );

    \I__5577\ : InMux
    port map (
            O => \N__31486\,
            I => \N__31428\
        );

    \I__5576\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31421\
        );

    \I__5575\ : InMux
    port map (
            O => \N__31484\,
            I => \N__31421\
        );

    \I__5574\ : InMux
    port map (
            O => \N__31483\,
            I => \N__31421\
        );

    \I__5573\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31410\
        );

    \I__5572\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31410\
        );

    \I__5571\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31410\
        );

    \I__5570\ : InMux
    port map (
            O => \N__31479\,
            I => \N__31410\
        );

    \I__5569\ : InMux
    port map (
            O => \N__31478\,
            I => \N__31410\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__31467\,
            I => \N__31405\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__31456\,
            I => \N__31405\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__31441\,
            I => \N__31402\
        );

    \I__5565\ : CascadeMux
    port map (
            O => \N__31440\,
            I => \N__31397\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__31437\,
            I => \N__31384\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__31428\,
            I => \N__31384\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__31421\,
            I => \N__31379\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__31410\,
            I => \N__31379\
        );

    \I__5560\ : Span4Mux_v
    port map (
            O => \N__31405\,
            I => \N__31374\
        );

    \I__5559\ : Span4Mux_v
    port map (
            O => \N__31402\,
            I => \N__31374\
        );

    \I__5558\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31371\
        );

    \I__5557\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31358\
        );

    \I__5556\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31358\
        );

    \I__5555\ : InMux
    port map (
            O => \N__31396\,
            I => \N__31358\
        );

    \I__5554\ : InMux
    port map (
            O => \N__31395\,
            I => \N__31358\
        );

    \I__5553\ : InMux
    port map (
            O => \N__31394\,
            I => \N__31358\
        );

    \I__5552\ : InMux
    port map (
            O => \N__31393\,
            I => \N__31358\
        );

    \I__5551\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31349\
        );

    \I__5550\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31349\
        );

    \I__5549\ : InMux
    port map (
            O => \N__31390\,
            I => \N__31349\
        );

    \I__5548\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31349\
        );

    \I__5547\ : Span4Mux_v
    port map (
            O => \N__31384\,
            I => \N__31346\
        );

    \I__5546\ : Span4Mux_v
    port map (
            O => \N__31379\,
            I => \N__31343\
        );

    \I__5545\ : Sp12to4
    port map (
            O => \N__31374\,
            I => \N__31340\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__31371\,
            I => measured_delay_hc_31
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__31358\,
            I => measured_delay_hc_31
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__31349\,
            I => measured_delay_hc_31
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__31346\,
            I => measured_delay_hc_31
        );

    \I__5540\ : Odrv4
    port map (
            O => \N__31343\,
            I => measured_delay_hc_31
        );

    \I__5539\ : Odrv12
    port map (
            O => \N__31340\,
            I => measured_delay_hc_31
        );

    \I__5538\ : InMux
    port map (
            O => \N__31327\,
            I => \N__31322\
        );

    \I__5537\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31319\
        );

    \I__5536\ : InMux
    port map (
            O => \N__31325\,
            I => \N__31314\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__31322\,
            I => \N__31311\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__31319\,
            I => \N__31308\
        );

    \I__5533\ : InMux
    port map (
            O => \N__31318\,
            I => \N__31305\
        );

    \I__5532\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31302\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__31314\,
            I => \N__31299\
        );

    \I__5530\ : Span4Mux_v
    port map (
            O => \N__31311\,
            I => \N__31294\
        );

    \I__5529\ : Span4Mux_h
    port map (
            O => \N__31308\,
            I => \N__31294\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__31305\,
            I => \N__31291\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__31302\,
            I => measured_delay_hc_3
        );

    \I__5526\ : Odrv4
    port map (
            O => \N__31299\,
            I => measured_delay_hc_3
        );

    \I__5525\ : Odrv4
    port map (
            O => \N__31294\,
            I => measured_delay_hc_3
        );

    \I__5524\ : Odrv12
    port map (
            O => \N__31291\,
            I => measured_delay_hc_3
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__31282\,
            I => \N__31275\
        );

    \I__5522\ : InMux
    port map (
            O => \N__31281\,
            I => \N__31272\
        );

    \I__5521\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31269\
        );

    \I__5520\ : InMux
    port map (
            O => \N__31279\,
            I => \N__31264\
        );

    \I__5519\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31264\
        );

    \I__5518\ : InMux
    port map (
            O => \N__31275\,
            I => \N__31261\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__31272\,
            I => \N__31258\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__31269\,
            I => \N__31253\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__31264\,
            I => \N__31253\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__31261\,
            I => measured_delay_hc_12
        );

    \I__5513\ : Odrv12
    port map (
            O => \N__31258\,
            I => measured_delay_hc_12
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__31253\,
            I => measured_delay_hc_12
        );

    \I__5511\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31241\
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__31245\,
            I => \N__31236\
        );

    \I__5509\ : InMux
    port map (
            O => \N__31244\,
            I => \N__31233\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__31241\,
            I => \N__31230\
        );

    \I__5507\ : InMux
    port map (
            O => \N__31240\,
            I => \N__31225\
        );

    \I__5506\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31225\
        );

    \I__5505\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31222\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__31233\,
            I => \N__31219\
        );

    \I__5503\ : Span4Mux_h
    port map (
            O => \N__31230\,
            I => \N__31216\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__31225\,
            I => \N__31213\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__31222\,
            I => measured_delay_hc_18
        );

    \I__5500\ : Odrv4
    port map (
            O => \N__31219\,
            I => measured_delay_hc_18
        );

    \I__5499\ : Odrv4
    port map (
            O => \N__31216\,
            I => measured_delay_hc_18
        );

    \I__5498\ : Odrv12
    port map (
            O => \N__31213\,
            I => measured_delay_hc_18
        );

    \I__5497\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31198\
        );

    \I__5496\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31192\
        );

    \I__5495\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31192\
        );

    \I__5494\ : CascadeMux
    port map (
            O => \N__31201\,
            I => \N__31189\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__31198\,
            I => \N__31186\
        );

    \I__5492\ : InMux
    port map (
            O => \N__31197\,
            I => \N__31183\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__31192\,
            I => \N__31180\
        );

    \I__5490\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31177\
        );

    \I__5489\ : Span4Mux_v
    port map (
            O => \N__31186\,
            I => \N__31170\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31170\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__31180\,
            I => \N__31170\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__31177\,
            I => measured_delay_hc_17
        );

    \I__5485\ : Odrv4
    port map (
            O => \N__31170\,
            I => measured_delay_hc_17
        );

    \I__5484\ : InMux
    port map (
            O => \N__31165\,
            I => \N__31160\
        );

    \I__5483\ : InMux
    port map (
            O => \N__31164\,
            I => \N__31157\
        );

    \I__5482\ : CascadeMux
    port map (
            O => \N__31163\,
            I => \N__31153\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__31160\,
            I => \N__31147\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__31157\,
            I => \N__31147\
        );

    \I__5479\ : InMux
    port map (
            O => \N__31156\,
            I => \N__31144\
        );

    \I__5478\ : InMux
    port map (
            O => \N__31153\,
            I => \N__31141\
        );

    \I__5477\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31138\
        );

    \I__5476\ : Span4Mux_h
    port map (
            O => \N__31147\,
            I => \N__31135\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__31144\,
            I => \N__31130\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__31141\,
            I => \N__31130\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__31138\,
            I => measured_delay_hc_5
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__31135\,
            I => measured_delay_hc_5
        );

    \I__5471\ : Odrv12
    port map (
            O => \N__31130\,
            I => measured_delay_hc_5
        );

    \I__5470\ : CascadeMux
    port map (
            O => \N__31123\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt9_0_cascade_\
        );

    \I__5469\ : InMux
    port map (
            O => \N__31120\,
            I => \N__31117\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__31117\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt15\
        );

    \I__5467\ : InMux
    port map (
            O => \N__31114\,
            I => \N__31111\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__31111\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1\
        );

    \I__5465\ : CascadeMux
    port map (
            O => \N__31108\,
            I => \N__31090\
        );

    \I__5464\ : CascadeMux
    port map (
            O => \N__31107\,
            I => \N__31087\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__31106\,
            I => \N__31084\
        );

    \I__5462\ : CascadeMux
    port map (
            O => \N__31105\,
            I => \N__31081\
        );

    \I__5461\ : CascadeMux
    port map (
            O => \N__31104\,
            I => \N__31074\
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__31103\,
            I => \N__31071\
        );

    \I__5459\ : CascadeMux
    port map (
            O => \N__31102\,
            I => \N__31068\
        );

    \I__5458\ : CascadeMux
    port map (
            O => \N__31101\,
            I => \N__31065\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__31100\,
            I => \N__31062\
        );

    \I__5456\ : CascadeMux
    port map (
            O => \N__31099\,
            I => \N__31059\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__31098\,
            I => \N__31056\
        );

    \I__5454\ : CascadeMux
    port map (
            O => \N__31097\,
            I => \N__31053\
        );

    \I__5453\ : CascadeMux
    port map (
            O => \N__31096\,
            I => \N__31050\
        );

    \I__5452\ : CascadeMux
    port map (
            O => \N__31095\,
            I => \N__31047\
        );

    \I__5451\ : CascadeMux
    port map (
            O => \N__31094\,
            I => \N__31044\
        );

    \I__5450\ : InMux
    port map (
            O => \N__31093\,
            I => \N__31027\
        );

    \I__5449\ : InMux
    port map (
            O => \N__31090\,
            I => \N__31027\
        );

    \I__5448\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31027\
        );

    \I__5447\ : InMux
    port map (
            O => \N__31084\,
            I => \N__31027\
        );

    \I__5446\ : InMux
    port map (
            O => \N__31081\,
            I => \N__31027\
        );

    \I__5445\ : InMux
    port map (
            O => \N__31080\,
            I => \N__31027\
        );

    \I__5444\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31027\
        );

    \I__5443\ : InMux
    port map (
            O => \N__31078\,
            I => \N__31027\
        );

    \I__5442\ : CascadeMux
    port map (
            O => \N__31077\,
            I => \N__31023\
        );

    \I__5441\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31013\
        );

    \I__5440\ : InMux
    port map (
            O => \N__31071\,
            I => \N__31013\
        );

    \I__5439\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31013\
        );

    \I__5438\ : InMux
    port map (
            O => \N__31065\,
            I => \N__31013\
        );

    \I__5437\ : InMux
    port map (
            O => \N__31062\,
            I => \N__31004\
        );

    \I__5436\ : InMux
    port map (
            O => \N__31059\,
            I => \N__31004\
        );

    \I__5435\ : InMux
    port map (
            O => \N__31056\,
            I => \N__31004\
        );

    \I__5434\ : InMux
    port map (
            O => \N__31053\,
            I => \N__31004\
        );

    \I__5433\ : InMux
    port map (
            O => \N__31050\,
            I => \N__30999\
        );

    \I__5432\ : InMux
    port map (
            O => \N__31047\,
            I => \N__30999\
        );

    \I__5431\ : InMux
    port map (
            O => \N__31044\,
            I => \N__30996\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__31027\,
            I => \N__30993\
        );

    \I__5429\ : InMux
    port map (
            O => \N__31026\,
            I => \N__30990\
        );

    \I__5428\ : InMux
    port map (
            O => \N__31023\,
            I => \N__30984\
        );

    \I__5427\ : InMux
    port map (
            O => \N__31022\,
            I => \N__30984\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__31013\,
            I => \N__30979\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__31004\,
            I => \N__30979\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__30999\,
            I => \N__30976\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__30996\,
            I => \N__30973\
        );

    \I__5422\ : Span4Mux_h
    port map (
            O => \N__30993\,
            I => \N__30967\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__30990\,
            I => \N__30967\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__30989\,
            I => \N__30964\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__30984\,
            I => \N__30959\
        );

    \I__5418\ : Span4Mux_v
    port map (
            O => \N__30979\,
            I => \N__30959\
        );

    \I__5417\ : Span4Mux_h
    port map (
            O => \N__30976\,
            I => \N__30954\
        );

    \I__5416\ : Span4Mux_h
    port map (
            O => \N__30973\,
            I => \N__30954\
        );

    \I__5415\ : InMux
    port map (
            O => \N__30972\,
            I => \N__30951\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__30967\,
            I => \N__30948\
        );

    \I__5413\ : InMux
    port map (
            O => \N__30964\,
            I => \N__30945\
        );

    \I__5412\ : Span4Mux_v
    port map (
            O => \N__30959\,
            I => \N__30942\
        );

    \I__5411\ : Sp12to4
    port map (
            O => \N__30954\,
            I => \N__30937\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__30951\,
            I => \N__30937\
        );

    \I__5409\ : Span4Mux_h
    port map (
            O => \N__30948\,
            I => \N__30934\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__30945\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__30942\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5406\ : Odrv12
    port map (
            O => \N__30937\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5405\ : Odrv4
    port map (
            O => \N__30934\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__30925\,
            I => \N__30919\
        );

    \I__5403\ : CascadeMux
    port map (
            O => \N__30924\,
            I => \N__30916\
        );

    \I__5402\ : CascadeMux
    port map (
            O => \N__30923\,
            I => \N__30913\
        );

    \I__5401\ : CascadeMux
    port map (
            O => \N__30922\,
            I => \N__30910\
        );

    \I__5400\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30883\
        );

    \I__5399\ : InMux
    port map (
            O => \N__30916\,
            I => \N__30883\
        );

    \I__5398\ : InMux
    port map (
            O => \N__30913\,
            I => \N__30883\
        );

    \I__5397\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30883\
        );

    \I__5396\ : InMux
    port map (
            O => \N__30909\,
            I => \N__30880\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30908\,
            I => \N__30863\
        );

    \I__5394\ : InMux
    port map (
            O => \N__30907\,
            I => \N__30863\
        );

    \I__5393\ : InMux
    port map (
            O => \N__30906\,
            I => \N__30863\
        );

    \I__5392\ : InMux
    port map (
            O => \N__30905\,
            I => \N__30863\
        );

    \I__5391\ : InMux
    port map (
            O => \N__30904\,
            I => \N__30863\
        );

    \I__5390\ : InMux
    port map (
            O => \N__30903\,
            I => \N__30863\
        );

    \I__5389\ : InMux
    port map (
            O => \N__30902\,
            I => \N__30863\
        );

    \I__5388\ : InMux
    port map (
            O => \N__30901\,
            I => \N__30863\
        );

    \I__5387\ : InMux
    port map (
            O => \N__30900\,
            I => \N__30854\
        );

    \I__5386\ : InMux
    port map (
            O => \N__30899\,
            I => \N__30854\
        );

    \I__5385\ : InMux
    port map (
            O => \N__30898\,
            I => \N__30854\
        );

    \I__5384\ : InMux
    port map (
            O => \N__30897\,
            I => \N__30854\
        );

    \I__5383\ : InMux
    port map (
            O => \N__30896\,
            I => \N__30851\
        );

    \I__5382\ : InMux
    port map (
            O => \N__30895\,
            I => \N__30848\
        );

    \I__5381\ : InMux
    port map (
            O => \N__30894\,
            I => \N__30845\
        );

    \I__5380\ : InMux
    port map (
            O => \N__30893\,
            I => \N__30838\
        );

    \I__5379\ : InMux
    port map (
            O => \N__30892\,
            I => \N__30838\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__30883\,
            I => \N__30829\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__30880\,
            I => \N__30829\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__30863\,
            I => \N__30829\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__30854\,
            I => \N__30829\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__30851\,
            I => \N__30826\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__30848\,
            I => \N__30821\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__30845\,
            I => \N__30821\
        );

    \I__5371\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30816\
        );

    \I__5370\ : InMux
    port map (
            O => \N__30843\,
            I => \N__30816\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30811\
        );

    \I__5368\ : Span4Mux_v
    port map (
            O => \N__30829\,
            I => \N__30811\
        );

    \I__5367\ : Span4Mux_v
    port map (
            O => \N__30826\,
            I => \N__30806\
        );

    \I__5366\ : Span4Mux_v
    port map (
            O => \N__30821\,
            I => \N__30806\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__30816\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__5364\ : Odrv4
    port map (
            O => \N__30811\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__5363\ : Odrv4
    port map (
            O => \N__30806\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__5362\ : InMux
    port map (
            O => \N__30799\,
            I => \N__30788\
        );

    \I__5361\ : InMux
    port map (
            O => \N__30798\,
            I => \N__30771\
        );

    \I__5360\ : InMux
    port map (
            O => \N__30797\,
            I => \N__30771\
        );

    \I__5359\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30771\
        );

    \I__5358\ : InMux
    port map (
            O => \N__30795\,
            I => \N__30771\
        );

    \I__5357\ : InMux
    port map (
            O => \N__30794\,
            I => \N__30771\
        );

    \I__5356\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30771\
        );

    \I__5355\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30771\
        );

    \I__5354\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30771\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__30788\,
            I => \N__30752\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__30771\,
            I => \N__30752\
        );

    \I__5351\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30749\
        );

    \I__5350\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30746\
        );

    \I__5349\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30741\
        );

    \I__5348\ : InMux
    port map (
            O => \N__30767\,
            I => \N__30741\
        );

    \I__5347\ : InMux
    port map (
            O => \N__30766\,
            I => \N__30724\
        );

    \I__5346\ : InMux
    port map (
            O => \N__30765\,
            I => \N__30724\
        );

    \I__5345\ : InMux
    port map (
            O => \N__30764\,
            I => \N__30724\
        );

    \I__5344\ : InMux
    port map (
            O => \N__30763\,
            I => \N__30724\
        );

    \I__5343\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30724\
        );

    \I__5342\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30724\
        );

    \I__5341\ : InMux
    port map (
            O => \N__30760\,
            I => \N__30724\
        );

    \I__5340\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30724\
        );

    \I__5339\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30721\
        );

    \I__5338\ : CascadeMux
    port map (
            O => \N__30757\,
            I => \N__30718\
        );

    \I__5337\ : Span4Mux_v
    port map (
            O => \N__30752\,
            I => \N__30712\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__30749\,
            I => \N__30712\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__30746\,
            I => \N__30709\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__30741\,
            I => \N__30702\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__30724\,
            I => \N__30702\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__30721\,
            I => \N__30702\
        );

    \I__5331\ : InMux
    port map (
            O => \N__30718\,
            I => \N__30697\
        );

    \I__5330\ : InMux
    port map (
            O => \N__30717\,
            I => \N__30697\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__30712\,
            I => \N__30692\
        );

    \I__5328\ : Span4Mux_v
    port map (
            O => \N__30709\,
            I => \N__30692\
        );

    \I__5327\ : Span4Mux_v
    port map (
            O => \N__30702\,
            I => \N__30689\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__30697\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5325\ : Odrv4
    port map (
            O => \N__30692\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__30689\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5323\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30678\
        );

    \I__5322\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30675\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__30678\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__30675\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0\
        );

    \I__5319\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30667\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30667\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__30664\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\
        );

    \I__5316\ : InMux
    port map (
            O => \N__30661\,
            I => \N__30658\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__30658\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12\
        );

    \I__5314\ : CascadeMux
    port map (
            O => \N__30655\,
            I => \N__30652\
        );

    \I__5313\ : InMux
    port map (
            O => \N__30652\,
            I => \N__30649\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__30649\,
            I => \N__30646\
        );

    \I__5311\ : Span4Mux_h
    port map (
            O => \N__30646\,
            I => \N__30643\
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__30643\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__30640\,
            I => \N__30637\
        );

    \I__5308\ : InMux
    port map (
            O => \N__30637\,
            I => \N__30634\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__30634\,
            I => \N__30631\
        );

    \I__5306\ : Odrv4
    port map (
            O => \N__30631\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__30628\,
            I => \N__30625\
        );

    \I__5304\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30622\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__30622\,
            I => \N__30619\
        );

    \I__5302\ : Span4Mux_h
    port map (
            O => \N__30619\,
            I => \N__30616\
        );

    \I__5301\ : Odrv4
    port map (
            O => \N__30616\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__5300\ : CEMux
    port map (
            O => \N__30613\,
            I => \N__30608\
        );

    \I__5299\ : CEMux
    port map (
            O => \N__30612\,
            I => \N__30605\
        );

    \I__5298\ : CEMux
    port map (
            O => \N__30611\,
            I => \N__30602\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__30608\,
            I => \N__30599\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__30605\,
            I => \N__30596\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__30602\,
            I => \N__30592\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__30599\,
            I => \N__30589\
        );

    \I__5293\ : Span4Mux_h
    port map (
            O => \N__30596\,
            I => \N__30586\
        );

    \I__5292\ : CEMux
    port map (
            O => \N__30595\,
            I => \N__30583\
        );

    \I__5291\ : Span4Mux_v
    port map (
            O => \N__30592\,
            I => \N__30580\
        );

    \I__5290\ : Span4Mux_h
    port map (
            O => \N__30589\,
            I => \N__30577\
        );

    \I__5289\ : Span4Mux_h
    port map (
            O => \N__30586\,
            I => \N__30574\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__30583\,
            I => \N__30571\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__30580\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5286\ : Odrv4
    port map (
            O => \N__30577\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__30574\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5284\ : Odrv12
    port map (
            O => \N__30571\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5283\ : CascadeMux
    port map (
            O => \N__30562\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_\
        );

    \I__5282\ : CascadeMux
    port map (
            O => \N__30559\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7_cascade_\
        );

    \I__5281\ : CascadeMux
    port map (
            O => \N__30556\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_\
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__30553\,
            I => \N__30546\
        );

    \I__5279\ : InMux
    port map (
            O => \N__30552\,
            I => \N__30540\
        );

    \I__5278\ : InMux
    port map (
            O => \N__30551\,
            I => \N__30533\
        );

    \I__5277\ : InMux
    port map (
            O => \N__30550\,
            I => \N__30533\
        );

    \I__5276\ : InMux
    port map (
            O => \N__30549\,
            I => \N__30533\
        );

    \I__5275\ : InMux
    port map (
            O => \N__30546\,
            I => \N__30530\
        );

    \I__5274\ : InMux
    port map (
            O => \N__30545\,
            I => \N__30523\
        );

    \I__5273\ : InMux
    port map (
            O => \N__30544\,
            I => \N__30523\
        );

    \I__5272\ : InMux
    port map (
            O => \N__30543\,
            I => \N__30523\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30520\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__30533\,
            I => \N__30517\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__30530\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__30523\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__5267\ : Odrv4
    port map (
            O => \N__30520\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__5266\ : Odrv12
    port map (
            O => \N__30517\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__5265\ : InMux
    port map (
            O => \N__30508\,
            I => \N__30505\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__30505\,
            I => \N__30502\
        );

    \I__5263\ : Span4Mux_h
    port map (
            O => \N__30502\,
            I => \N__30499\
        );

    \I__5262\ : Span4Mux_v
    port map (
            O => \N__30499\,
            I => \N__30493\
        );

    \I__5261\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30490\
        );

    \I__5260\ : InMux
    port map (
            O => \N__30497\,
            I => \N__30487\
        );

    \I__5259\ : InMux
    port map (
            O => \N__30496\,
            I => \N__30484\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__30493\,
            I => \N__30481\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__30490\,
            I => \N__30478\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__30487\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__30484\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__30481\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__30478\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5252\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30466\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__30466\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3\
        );

    \I__5250\ : CascadeMux
    port map (
            O => \N__30463\,
            I => \N__30460\
        );

    \I__5249\ : InMux
    port map (
            O => \N__30460\,
            I => \N__30457\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__30457\,
            I => \N__30454\
        );

    \I__5247\ : Span4Mux_h
    port map (
            O => \N__30454\,
            I => \N__30451\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__30451\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__5245\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30430\
        );

    \I__5244\ : InMux
    port map (
            O => \N__30447\,
            I => \N__30430\
        );

    \I__5243\ : InMux
    port map (
            O => \N__30446\,
            I => \N__30405\
        );

    \I__5242\ : InMux
    port map (
            O => \N__30445\,
            I => \N__30405\
        );

    \I__5241\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30405\
        );

    \I__5240\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30405\
        );

    \I__5239\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30405\
        );

    \I__5238\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30405\
        );

    \I__5237\ : InMux
    port map (
            O => \N__30440\,
            I => \N__30405\
        );

    \I__5236\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30405\
        );

    \I__5235\ : InMux
    port map (
            O => \N__30438\,
            I => \N__30402\
        );

    \I__5234\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30397\
        );

    \I__5233\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30397\
        );

    \I__5232\ : InMux
    port map (
            O => \N__30435\,
            I => \N__30394\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__30430\,
            I => \N__30391\
        );

    \I__5230\ : InMux
    port map (
            O => \N__30429\,
            I => \N__30372\
        );

    \I__5229\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30372\
        );

    \I__5228\ : InMux
    port map (
            O => \N__30427\,
            I => \N__30372\
        );

    \I__5227\ : InMux
    port map (
            O => \N__30426\,
            I => \N__30372\
        );

    \I__5226\ : InMux
    port map (
            O => \N__30425\,
            I => \N__30372\
        );

    \I__5225\ : InMux
    port map (
            O => \N__30424\,
            I => \N__30372\
        );

    \I__5224\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30372\
        );

    \I__5223\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30372\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__30405\,
            I => \N__30369\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__30402\,
            I => \N__30366\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__30397\,
            I => \N__30361\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__30394\,
            I => \N__30361\
        );

    \I__5218\ : Span4Mux_v
    port map (
            O => \N__30391\,
            I => \N__30358\
        );

    \I__5217\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30353\
        );

    \I__5216\ : InMux
    port map (
            O => \N__30389\,
            I => \N__30353\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__30372\,
            I => \N__30346\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__30369\,
            I => \N__30346\
        );

    \I__5213\ : Span4Mux_h
    port map (
            O => \N__30366\,
            I => \N__30346\
        );

    \I__5212\ : Sp12to4
    port map (
            O => \N__30361\,
            I => \N__30343\
        );

    \I__5211\ : Span4Mux_h
    port map (
            O => \N__30358\,
            I => \N__30340\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__30353\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__30346\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5208\ : Odrv12
    port map (
            O => \N__30343\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5207\ : Odrv4
    port map (
            O => \N__30340\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__5206\ : CascadeMux
    port map (
            O => \N__30331\,
            I => \N__30328\
        );

    \I__5205\ : InMux
    port map (
            O => \N__30328\,
            I => \N__30310\
        );

    \I__5204\ : InMux
    port map (
            O => \N__30327\,
            I => \N__30310\
        );

    \I__5203\ : CascadeMux
    port map (
            O => \N__30326\,
            I => \N__30304\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__30325\,
            I => \N__30301\
        );

    \I__5201\ : CascadeMux
    port map (
            O => \N__30324\,
            I => \N__30298\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__30323\,
            I => \N__30295\
        );

    \I__5199\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30274\
        );

    \I__5198\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30274\
        );

    \I__5197\ : InMux
    port map (
            O => \N__30320\,
            I => \N__30274\
        );

    \I__5196\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30274\
        );

    \I__5195\ : InMux
    port map (
            O => \N__30318\,
            I => \N__30274\
        );

    \I__5194\ : InMux
    port map (
            O => \N__30317\,
            I => \N__30274\
        );

    \I__5193\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30274\
        );

    \I__5192\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30274\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__30310\,
            I => \N__30271\
        );

    \I__5190\ : InMux
    port map (
            O => \N__30309\,
            I => \N__30268\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__30308\,
            I => \N__30265\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__30307\,
            I => \N__30262\
        );

    \I__5187\ : InMux
    port map (
            O => \N__30304\,
            I => \N__30243\
        );

    \I__5186\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30243\
        );

    \I__5185\ : InMux
    port map (
            O => \N__30298\,
            I => \N__30243\
        );

    \I__5184\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30243\
        );

    \I__5183\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30243\
        );

    \I__5182\ : InMux
    port map (
            O => \N__30293\,
            I => \N__30243\
        );

    \I__5181\ : InMux
    port map (
            O => \N__30292\,
            I => \N__30243\
        );

    \I__5180\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30243\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__30274\,
            I => \N__30240\
        );

    \I__5178\ : Span4Mux_v
    port map (
            O => \N__30271\,
            I => \N__30234\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__30268\,
            I => \N__30234\
        );

    \I__5176\ : InMux
    port map (
            O => \N__30265\,
            I => \N__30229\
        );

    \I__5175\ : InMux
    port map (
            O => \N__30262\,
            I => \N__30229\
        );

    \I__5174\ : InMux
    port map (
            O => \N__30261\,
            I => \N__30224\
        );

    \I__5173\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30224\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__30243\,
            I => \N__30221\
        );

    \I__5171\ : Span4Mux_v
    port map (
            O => \N__30240\,
            I => \N__30218\
        );

    \I__5170\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30215\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__30234\,
            I => \N__30212\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__30229\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__30224\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__30221\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5165\ : Odrv4
    port map (
            O => \N__30218\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__30215\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5163\ : Odrv4
    port map (
            O => \N__30212\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__5162\ : CascadeMux
    port map (
            O => \N__30199\,
            I => \N__30176\
        );

    \I__5161\ : CascadeMux
    port map (
            O => \N__30198\,
            I => \N__30173\
        );

    \I__5160\ : CascadeMux
    port map (
            O => \N__30197\,
            I => \N__30170\
        );

    \I__5159\ : CascadeMux
    port map (
            O => \N__30196\,
            I => \N__30167\
        );

    \I__5158\ : InMux
    port map (
            O => \N__30195\,
            I => \N__30149\
        );

    \I__5157\ : InMux
    port map (
            O => \N__30194\,
            I => \N__30149\
        );

    \I__5156\ : InMux
    port map (
            O => \N__30193\,
            I => \N__30149\
        );

    \I__5155\ : InMux
    port map (
            O => \N__30192\,
            I => \N__30149\
        );

    \I__5154\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30149\
        );

    \I__5153\ : InMux
    port map (
            O => \N__30190\,
            I => \N__30149\
        );

    \I__5152\ : InMux
    port map (
            O => \N__30189\,
            I => \N__30149\
        );

    \I__5151\ : InMux
    port map (
            O => \N__30188\,
            I => \N__30149\
        );

    \I__5150\ : InMux
    port map (
            O => \N__30187\,
            I => \N__30143\
        );

    \I__5149\ : InMux
    port map (
            O => \N__30186\,
            I => \N__30143\
        );

    \I__5148\ : CascadeMux
    port map (
            O => \N__30185\,
            I => \N__30140\
        );

    \I__5147\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30134\
        );

    \I__5146\ : InMux
    port map (
            O => \N__30183\,
            I => \N__30134\
        );

    \I__5145\ : InMux
    port map (
            O => \N__30182\,
            I => \N__30117\
        );

    \I__5144\ : InMux
    port map (
            O => \N__30181\,
            I => \N__30117\
        );

    \I__5143\ : InMux
    port map (
            O => \N__30180\,
            I => \N__30117\
        );

    \I__5142\ : InMux
    port map (
            O => \N__30179\,
            I => \N__30117\
        );

    \I__5141\ : InMux
    port map (
            O => \N__30176\,
            I => \N__30117\
        );

    \I__5140\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30117\
        );

    \I__5139\ : InMux
    port map (
            O => \N__30170\,
            I => \N__30117\
        );

    \I__5138\ : InMux
    port map (
            O => \N__30167\,
            I => \N__30117\
        );

    \I__5137\ : InMux
    port map (
            O => \N__30166\,
            I => \N__30114\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__30149\,
            I => \N__30111\
        );

    \I__5135\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30108\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__30143\,
            I => \N__30105\
        );

    \I__5133\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30100\
        );

    \I__5132\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30100\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__30134\,
            I => \N__30097\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__30117\,
            I => \N__30092\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__30114\,
            I => \N__30092\
        );

    \I__5128\ : Span4Mux_v
    port map (
            O => \N__30111\,
            I => \N__30085\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__30108\,
            I => \N__30085\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__30105\,
            I => \N__30085\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__30100\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__5124\ : Odrv12
    port map (
            O => \N__30097\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__30092\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__30085\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__5121\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30072\
        );

    \I__5120\ : InMux
    port map (
            O => \N__30075\,
            I => \N__30069\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__30072\,
            I => \N__30066\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__30069\,
            I => \N__30062\
        );

    \I__5117\ : Span12Mux_h
    port map (
            O => \N__30066\,
            I => \N__30058\
        );

    \I__5116\ : InMux
    port map (
            O => \N__30065\,
            I => \N__30055\
        );

    \I__5115\ : Span4Mux_v
    port map (
            O => \N__30062\,
            I => \N__30052\
        );

    \I__5114\ : InMux
    port map (
            O => \N__30061\,
            I => \N__30049\
        );

    \I__5113\ : Odrv12
    port map (
            O => \N__30058\,
            I => \phase_controller_inst2.stoper_hc.time_passed11\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__30055\,
            I => \phase_controller_inst2.stoper_hc.time_passed11\
        );

    \I__5111\ : Odrv4
    port map (
            O => \N__30052\,
            I => \phase_controller_inst2.stoper_hc.time_passed11\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__30049\,
            I => \phase_controller_inst2.stoper_hc.time_passed11\
        );

    \I__5109\ : InMux
    port map (
            O => \N__30040\,
            I => \N__30037\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__30037\,
            I => \N__30034\
        );

    \I__5107\ : Span4Mux_v
    port map (
            O => \N__30034\,
            I => \N__30028\
        );

    \I__5106\ : InMux
    port map (
            O => \N__30033\,
            I => \N__30021\
        );

    \I__5105\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30021\
        );

    \I__5104\ : InMux
    port map (
            O => \N__30031\,
            I => \N__30021\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__30028\,
            I => \N__30016\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__30021\,
            I => \N__30013\
        );

    \I__5101\ : InMux
    port map (
            O => \N__30020\,
            I => \N__30008\
        );

    \I__5100\ : InMux
    port map (
            O => \N__30019\,
            I => \N__30008\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__30016\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__30013\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__30008\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5096\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29998\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__29998\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0\
        );

    \I__5094\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29984\
        );

    \I__5093\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29984\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__29993\,
            I => \N__29978\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__29992\,
            I => \N__29975\
        );

    \I__5090\ : CascadeMux
    port map (
            O => \N__29991\,
            I => \N__29972\
        );

    \I__5089\ : CascadeMux
    port map (
            O => \N__29990\,
            I => \N__29969\
        );

    \I__5088\ : CascadeMux
    port map (
            O => \N__29989\,
            I => \N__29966\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__29984\,
            I => \N__29960\
        );

    \I__5086\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29942\
        );

    \I__5085\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29942\
        );

    \I__5084\ : InMux
    port map (
            O => \N__29981\,
            I => \N__29942\
        );

    \I__5083\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29942\
        );

    \I__5082\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29942\
        );

    \I__5081\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29942\
        );

    \I__5080\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29931\
        );

    \I__5079\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29931\
        );

    \I__5078\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29931\
        );

    \I__5077\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29931\
        );

    \I__5076\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29931\
        );

    \I__5075\ : Span4Mux_v
    port map (
            O => \N__29960\,
            I => \N__29928\
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__29959\,
            I => \N__29923\
        );

    \I__5073\ : CascadeMux
    port map (
            O => \N__29958\,
            I => \N__29920\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__29957\,
            I => \N__29917\
        );

    \I__5071\ : CascadeMux
    port map (
            O => \N__29956\,
            I => \N__29914\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__29955\,
            I => \N__29911\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__29942\,
            I => \N__29900\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__29931\,
            I => \N__29900\
        );

    \I__5067\ : Span4Mux_h
    port map (
            O => \N__29928\,
            I => \N__29900\
        );

    \I__5066\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29895\
        );

    \I__5065\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29895\
        );

    \I__5064\ : InMux
    port map (
            O => \N__29923\,
            I => \N__29892\
        );

    \I__5063\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29877\
        );

    \I__5062\ : InMux
    port map (
            O => \N__29917\,
            I => \N__29877\
        );

    \I__5061\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29877\
        );

    \I__5060\ : InMux
    port map (
            O => \N__29911\,
            I => \N__29877\
        );

    \I__5059\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29877\
        );

    \I__5058\ : InMux
    port map (
            O => \N__29909\,
            I => \N__29877\
        );

    \I__5057\ : InMux
    port map (
            O => \N__29908\,
            I => \N__29877\
        );

    \I__5056\ : InMux
    port map (
            O => \N__29907\,
            I => \N__29874\
        );

    \I__5055\ : Span4Mux_v
    port map (
            O => \N__29900\,
            I => \N__29869\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__29895\,
            I => \N__29869\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__29892\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__29877\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__29874\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5050\ : Odrv4
    port map (
            O => \N__29869\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5049\ : InMux
    port map (
            O => \N__29860\,
            I => \N__29855\
        );

    \I__5048\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29852\
        );

    \I__5047\ : InMux
    port map (
            O => \N__29858\,
            I => \N__29849\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__29855\,
            I => \N__29845\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__29852\,
            I => \N__29840\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__29849\,
            I => \N__29840\
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__29848\,
            I => \N__29837\
        );

    \I__5042\ : Span4Mux_v
    port map (
            O => \N__29845\,
            I => \N__29830\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__29840\,
            I => \N__29830\
        );

    \I__5040\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29827\
        );

    \I__5039\ : InMux
    port map (
            O => \N__29836\,
            I => \N__29822\
        );

    \I__5038\ : InMux
    port map (
            O => \N__29835\,
            I => \N__29822\
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__29830\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__29827\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__29822\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5034\ : InMux
    port map (
            O => \N__29815\,
            I => \N__29794\
        );

    \I__5033\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29779\
        );

    \I__5032\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29779\
        );

    \I__5031\ : InMux
    port map (
            O => \N__29812\,
            I => \N__29779\
        );

    \I__5030\ : InMux
    port map (
            O => \N__29811\,
            I => \N__29779\
        );

    \I__5029\ : InMux
    port map (
            O => \N__29810\,
            I => \N__29779\
        );

    \I__5028\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29779\
        );

    \I__5027\ : InMux
    port map (
            O => \N__29808\,
            I => \N__29779\
        );

    \I__5026\ : InMux
    port map (
            O => \N__29807\,
            I => \N__29766\
        );

    \I__5025\ : InMux
    port map (
            O => \N__29806\,
            I => \N__29766\
        );

    \I__5024\ : InMux
    port map (
            O => \N__29805\,
            I => \N__29766\
        );

    \I__5023\ : InMux
    port map (
            O => \N__29804\,
            I => \N__29766\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29803\,
            I => \N__29766\
        );

    \I__5021\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29766\
        );

    \I__5020\ : InMux
    port map (
            O => \N__29801\,
            I => \N__29755\
        );

    \I__5019\ : InMux
    port map (
            O => \N__29800\,
            I => \N__29755\
        );

    \I__5018\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29755\
        );

    \I__5017\ : InMux
    port map (
            O => \N__29798\,
            I => \N__29755\
        );

    \I__5016\ : InMux
    port map (
            O => \N__29797\,
            I => \N__29755\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__29794\,
            I => \N__29747\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__29779\,
            I => \N__29747\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__29766\,
            I => \N__29742\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__29755\,
            I => \N__29742\
        );

    \I__5011\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29735\
        );

    \I__5010\ : InMux
    port map (
            O => \N__29753\,
            I => \N__29735\
        );

    \I__5009\ : InMux
    port map (
            O => \N__29752\,
            I => \N__29735\
        );

    \I__5008\ : Span4Mux_v
    port map (
            O => \N__29747\,
            I => \N__29726\
        );

    \I__5007\ : Span4Mux_v
    port map (
            O => \N__29742\,
            I => \N__29726\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__29735\,
            I => \N__29726\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__29734\,
            I => \N__29723\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__29733\,
            I => \N__29720\
        );

    \I__5003\ : Span4Mux_h
    port map (
            O => \N__29726\,
            I => \N__29717\
        );

    \I__5002\ : InMux
    port map (
            O => \N__29723\,
            I => \N__29714\
        );

    \I__5001\ : InMux
    port map (
            O => \N__29720\,
            I => \N__29711\
        );

    \I__5000\ : Span4Mux_v
    port map (
            O => \N__29717\,
            I => \N__29708\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__29714\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__29711\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__29708\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__4996\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29686\
        );

    \I__4995\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29671\
        );

    \I__4994\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29671\
        );

    \I__4993\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29671\
        );

    \I__4992\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29671\
        );

    \I__4991\ : InMux
    port map (
            O => \N__29696\,
            I => \N__29671\
        );

    \I__4990\ : InMux
    port map (
            O => \N__29695\,
            I => \N__29671\
        );

    \I__4989\ : InMux
    port map (
            O => \N__29694\,
            I => \N__29671\
        );

    \I__4988\ : InMux
    port map (
            O => \N__29693\,
            I => \N__29660\
        );

    \I__4987\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29660\
        );

    \I__4986\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29660\
        );

    \I__4985\ : InMux
    port map (
            O => \N__29690\,
            I => \N__29660\
        );

    \I__4984\ : InMux
    port map (
            O => \N__29689\,
            I => \N__29660\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__29686\,
            I => \N__29646\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__29671\,
            I => \N__29646\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__29660\,
            I => \N__29643\
        );

    \I__4980\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29640\
        );

    \I__4979\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29635\
        );

    \I__4978\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29635\
        );

    \I__4977\ : InMux
    port map (
            O => \N__29656\,
            I => \N__29622\
        );

    \I__4976\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29622\
        );

    \I__4975\ : InMux
    port map (
            O => \N__29654\,
            I => \N__29622\
        );

    \I__4974\ : InMux
    port map (
            O => \N__29653\,
            I => \N__29622\
        );

    \I__4973\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29622\
        );

    \I__4972\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29622\
        );

    \I__4971\ : Span4Mux_v
    port map (
            O => \N__29646\,
            I => \N__29613\
        );

    \I__4970\ : Span4Mux_v
    port map (
            O => \N__29643\,
            I => \N__29613\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__29640\,
            I => \N__29613\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__29635\,
            I => \N__29613\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__29622\,
            I => \N__29608\
        );

    \I__4966\ : Span4Mux_h
    port map (
            O => \N__29613\,
            I => \N__29605\
        );

    \I__4965\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29600\
        );

    \I__4964\ : InMux
    port map (
            O => \N__29611\,
            I => \N__29600\
        );

    \I__4963\ : Span4Mux_h
    port map (
            O => \N__29608\,
            I => \N__29597\
        );

    \I__4962\ : Span4Mux_v
    port map (
            O => \N__29605\,
            I => \N__29594\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__29600\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__4960\ : Odrv4
    port map (
            O => \N__29597\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__4959\ : Odrv4
    port map (
            O => \N__29594\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__4958\ : CascadeMux
    port map (
            O => \N__29587\,
            I => \N__29584\
        );

    \I__4957\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29581\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__29581\,
            I => \N__29578\
        );

    \I__4955\ : Span4Mux_v
    port map (
            O => \N__29578\,
            I => \N__29575\
        );

    \I__4954\ : Odrv4
    port map (
            O => \N__29575\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__29572\,
            I => \N__29569\
        );

    \I__4952\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29566\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__29566\,
            I => \N__29563\
        );

    \I__4950\ : Span4Mux_h
    port map (
            O => \N__29563\,
            I => \N__29560\
        );

    \I__4949\ : Odrv4
    port map (
            O => \N__29560\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__4948\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29554\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__29554\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__4946\ : CascadeMux
    port map (
            O => \N__29551\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__29548\,
            I => \N__29545\
        );

    \I__4944\ : InMux
    port map (
            O => \N__29545\,
            I => \N__29542\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__29542\,
            I => \N__29539\
        );

    \I__4942\ : Odrv4
    port map (
            O => \N__29539\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__4941\ : CascadeMux
    port map (
            O => \N__29536\,
            I => \N__29533\
        );

    \I__4940\ : InMux
    port map (
            O => \N__29533\,
            I => \N__29530\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__29530\,
            I => \N__29527\
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__29527\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__4937\ : CascadeMux
    port map (
            O => \N__29524\,
            I => \N__29521\
        );

    \I__4936\ : InMux
    port map (
            O => \N__29521\,
            I => \N__29518\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__29518\,
            I => \N__29515\
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__29515\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__4933\ : CascadeMux
    port map (
            O => \N__29512\,
            I => \N__29509\
        );

    \I__4932\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29506\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__29506\,
            I => \N__29503\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__29503\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__4929\ : CascadeMux
    port map (
            O => \N__29500\,
            I => \delay_measurement_inst.N_265_cascade_\
        );

    \I__4928\ : InMux
    port map (
            O => \N__29497\,
            I => \N__29491\
        );

    \I__4927\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29491\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__29491\,
            I => \N__29484\
        );

    \I__4925\ : InMux
    port map (
            O => \N__29490\,
            I => \N__29475\
        );

    \I__4924\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29475\
        );

    \I__4923\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29475\
        );

    \I__4922\ : InMux
    port map (
            O => \N__29487\,
            I => \N__29475\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__29484\,
            I => \delay_measurement_inst.N_270\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__29475\,
            I => \delay_measurement_inst.N_270\
        );

    \I__4919\ : InMux
    port map (
            O => \N__29470\,
            I => \N__29467\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__29467\,
            I => \N__29464\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__29464\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\
        );

    \I__4916\ : InMux
    port map (
            O => \N__29461\,
            I => \N__29458\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__29458\,
            I => \N__29453\
        );

    \I__4914\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29450\
        );

    \I__4913\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29447\
        );

    \I__4912\ : Span4Mux_v
    port map (
            O => \N__29453\,
            I => \N__29444\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__29450\,
            I => \N__29440\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__29447\,
            I => \N__29437\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__29444\,
            I => \N__29434\
        );

    \I__4908\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29431\
        );

    \I__4907\ : Span4Mux_v
    port map (
            O => \N__29440\,
            I => \N__29426\
        );

    \I__4906\ : Span4Mux_v
    port map (
            O => \N__29437\,
            I => \N__29426\
        );

    \I__4905\ : Odrv4
    port map (
            O => \N__29434\,
            I => measured_delay_tr_17
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__29431\,
            I => measured_delay_tr_17
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__29426\,
            I => measured_delay_tr_17
        );

    \I__4902\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29414\
        );

    \I__4901\ : InMux
    port map (
            O => \N__29418\,
            I => \N__29411\
        );

    \I__4900\ : InMux
    port map (
            O => \N__29417\,
            I => \N__29408\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__29414\,
            I => \N__29404\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__29411\,
            I => \N__29399\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__29408\,
            I => \N__29399\
        );

    \I__4896\ : InMux
    port map (
            O => \N__29407\,
            I => \N__29396\
        );

    \I__4895\ : Span4Mux_h
    port map (
            O => \N__29404\,
            I => \N__29391\
        );

    \I__4894\ : Span4Mux_h
    port map (
            O => \N__29399\,
            I => \N__29391\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__29396\,
            I => measured_delay_tr_18
        );

    \I__4892\ : Odrv4
    port map (
            O => \N__29391\,
            I => measured_delay_tr_18
        );

    \I__4891\ : InMux
    port map (
            O => \N__29386\,
            I => \N__29376\
        );

    \I__4890\ : InMux
    port map (
            O => \N__29385\,
            I => \N__29376\
        );

    \I__4889\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29376\
        );

    \I__4888\ : InMux
    port map (
            O => \N__29383\,
            I => \N__29370\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__29376\,
            I => \N__29367\
        );

    \I__4886\ : InMux
    port map (
            O => \N__29375\,
            I => \N__29362\
        );

    \I__4885\ : InMux
    port map (
            O => \N__29374\,
            I => \N__29362\
        );

    \I__4884\ : InMux
    port map (
            O => \N__29373\,
            I => \N__29359\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__29370\,
            I => \N__29354\
        );

    \I__4882\ : Span4Mux_v
    port map (
            O => \N__29367\,
            I => \N__29347\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__29362\,
            I => \N__29347\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__29359\,
            I => \N__29347\
        );

    \I__4879\ : InMux
    port map (
            O => \N__29358\,
            I => \N__29342\
        );

    \I__4878\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29342\
        );

    \I__4877\ : Odrv4
    port map (
            O => \N__29354\,
            I => \delay_measurement_inst.N_325\
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__29347\,
            I => \delay_measurement_inst.N_325\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__29342\,
            I => \delay_measurement_inst.N_325\
        );

    \I__4874\ : CascadeMux
    port map (
            O => \N__29335\,
            I => \N__29330\
        );

    \I__4873\ : InMux
    port map (
            O => \N__29334\,
            I => \N__29326\
        );

    \I__4872\ : InMux
    port map (
            O => \N__29333\,
            I => \N__29323\
        );

    \I__4871\ : InMux
    port map (
            O => \N__29330\,
            I => \N__29320\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__29329\,
            I => \N__29317\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__29326\,
            I => \N__29314\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__29323\,
            I => \N__29309\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__29320\,
            I => \N__29309\
        );

    \I__4866\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29306\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__29314\,
            I => \N__29301\
        );

    \I__4864\ : Span4Mux_h
    port map (
            O => \N__29309\,
            I => \N__29301\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__29306\,
            I => measured_delay_tr_19
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__29301\,
            I => measured_delay_tr_19
        );

    \I__4861\ : CEMux
    port map (
            O => \N__29296\,
            I => \N__29293\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__29293\,
            I => \N__29290\
        );

    \I__4859\ : Sp12to4
    port map (
            O => \N__29290\,
            I => \N__29284\
        );

    \I__4858\ : CEMux
    port map (
            O => \N__29289\,
            I => \N__29281\
        );

    \I__4857\ : CEMux
    port map (
            O => \N__29288\,
            I => \N__29278\
        );

    \I__4856\ : CEMux
    port map (
            O => \N__29287\,
            I => \N__29275\
        );

    \I__4855\ : Odrv12
    port map (
            O => \N__29284\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__29281\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__29278\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__29275\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__4851\ : InMux
    port map (
            O => \N__29266\,
            I => \N__29263\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__29263\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__4849\ : CascadeMux
    port map (
            O => \N__29260\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_\
        );

    \I__4848\ : InMux
    port map (
            O => \N__29257\,
            I => \N__29254\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__29254\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5\
        );

    \I__4846\ : CascadeMux
    port map (
            O => \N__29251\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_\
        );

    \I__4845\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29244\
        );

    \I__4844\ : InMux
    port map (
            O => \N__29247\,
            I => \N__29241\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__29244\,
            I => \N__29236\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__29241\,
            I => \N__29236\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__29236\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i\
        );

    \I__4840\ : CascadeMux
    port map (
            O => \N__29233\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_\
        );

    \I__4839\ : InMux
    port map (
            O => \N__29230\,
            I => \N__29227\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__29227\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5\
        );

    \I__4837\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29218\
        );

    \I__4836\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29218\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__29218\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7\
        );

    \I__4834\ : InMux
    port map (
            O => \N__29215\,
            I => \N__29204\
        );

    \I__4833\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29204\
        );

    \I__4832\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29195\
        );

    \I__4831\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29195\
        );

    \I__4830\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29195\
        );

    \I__4829\ : InMux
    port map (
            O => \N__29210\,
            I => \N__29195\
        );

    \I__4828\ : InMux
    port map (
            O => \N__29209\,
            I => \N__29192\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__29204\,
            I => \delay_measurement_inst.N_299\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__29195\,
            I => \delay_measurement_inst.N_299\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__29192\,
            I => \delay_measurement_inst.N_299\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__29185\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\
        );

    \I__4823\ : InMux
    port map (
            O => \N__29182\,
            I => \N__29179\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__29179\,
            I => \delay_measurement_inst.delay_tr_timer.N_287_4\
        );

    \I__4821\ : InMux
    port map (
            O => \N__29176\,
            I => \N__29173\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__29173\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\
        );

    \I__4819\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29167\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__29167\,
            I => \N__29163\
        );

    \I__4817\ : InMux
    port map (
            O => \N__29166\,
            I => \N__29159\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__29163\,
            I => \N__29156\
        );

    \I__4815\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29153\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__29159\,
            I => \delay_measurement_inst.N_265\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__29156\,
            I => \delay_measurement_inst.N_265\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__29153\,
            I => \delay_measurement_inst.N_265\
        );

    \I__4811\ : InMux
    port map (
            O => \N__29146\,
            I => \N__29143\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__29143\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__4809\ : InMux
    port map (
            O => \N__29140\,
            I => \N__29137\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__29137\,
            I => \N__29134\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__29134\,
            I => \N__29131\
        );

    \I__4806\ : Odrv4
    port map (
            O => \N__29131\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__4805\ : InMux
    port map (
            O => \N__29128\,
            I => \N__29125\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__29125\,
            I => \N__29122\
        );

    \I__4803\ : Odrv4
    port map (
            O => \N__29122\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__29119\,
            I => \delay_measurement_inst.delay_tr_timer.N_287_4_cascade_\
        );

    \I__4801\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29113\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__29113\,
            I => \N__29110\
        );

    \I__4799\ : Odrv4
    port map (
            O => \N__29110\,
            I => \delay_measurement_inst.delay_tr_timer.N_290\
        );

    \I__4798\ : CascadeMux
    port map (
            O => \N__29107\,
            I => \N__29104\
        );

    \I__4797\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29101\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__29101\,
            I => \delay_measurement_inst.N_59\
        );

    \I__4795\ : InMux
    port map (
            O => \N__29098\,
            I => \N__29092\
        );

    \I__4794\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29092\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__29092\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\
        );

    \I__4792\ : CascadeMux
    port map (
            O => \N__29089\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\
        );

    \I__4791\ : InMux
    port map (
            O => \N__29086\,
            I => \N__29083\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__29083\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__4789\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29077\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__29077\,
            I => \N__29074\
        );

    \I__4787\ : Odrv12
    port map (
            O => \N__29074\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\
        );

    \I__4786\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29068\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29065\
        );

    \I__4784\ : Odrv12
    port map (
            O => \N__29065\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\
        );

    \I__4783\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29059\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__29059\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__29056\,
            I => \N__29048\
        );

    \I__4780\ : CascadeMux
    port map (
            O => \N__29055\,
            I => \N__29045\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__29054\,
            I => \N__29042\
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__29053\,
            I => \N__29039\
        );

    \I__4777\ : InMux
    port map (
            O => \N__29052\,
            I => \N__29030\
        );

    \I__4776\ : InMux
    port map (
            O => \N__29051\,
            I => \N__29030\
        );

    \I__4775\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29030\
        );

    \I__4774\ : InMux
    port map (
            O => \N__29045\,
            I => \N__29030\
        );

    \I__4773\ : InMux
    port map (
            O => \N__29042\,
            I => \N__29023\
        );

    \I__4772\ : InMux
    port map (
            O => \N__29039\,
            I => \N__29023\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__29030\,
            I => \N__29020\
        );

    \I__4770\ : InMux
    port map (
            O => \N__29029\,
            I => \N__29017\
        );

    \I__4769\ : InMux
    port map (
            O => \N__29028\,
            I => \N__29014\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__29023\,
            I => \N__29005\
        );

    \I__4767\ : Span4Mux_h
    port map (
            O => \N__29020\,
            I => \N__29005\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__29017\,
            I => \N__29005\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__29014\,
            I => \N__29005\
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__29005\,
            I => \delay_measurement_inst.N_267\
        );

    \I__4763\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__28999\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\
        );

    \I__4761\ : CascadeMux
    port map (
            O => \N__28996\,
            I => \N__28993\
        );

    \I__4760\ : InMux
    port map (
            O => \N__28993\,
            I => \N__28990\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__28990\,
            I => \N__28987\
        );

    \I__4758\ : Odrv4
    port map (
            O => \N__28987\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__4757\ : CascadeMux
    port map (
            O => \N__28984\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\
        );

    \I__4756\ : CascadeMux
    port map (
            O => \N__28981\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__28978\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__4754\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28972\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__28972\,
            I => \current_shift_inst.PI_CTRL.N_72\
        );

    \I__4752\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28966\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__28966\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__28963\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\
        );

    \I__4749\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28957\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__28957\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__28954\,
            I => \N__28951\
        );

    \I__4746\ : InMux
    port map (
            O => \N__28951\,
            I => \N__28948\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28948\,
            I => \N__28945\
        );

    \I__4744\ : Span4Mux_h
    port map (
            O => \N__28945\,
            I => \N__28942\
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__28942\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__28939\,
            I => \N__28936\
        );

    \I__4741\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28933\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__28933\,
            I => \N__28930\
        );

    \I__4739\ : Span4Mux_h
    port map (
            O => \N__28930\,
            I => \N__28927\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__28927\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__28924\,
            I => \N__28921\
        );

    \I__4736\ : InMux
    port map (
            O => \N__28921\,
            I => \N__28918\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__28918\,
            I => \N__28915\
        );

    \I__4734\ : Span4Mux_h
    port map (
            O => \N__28915\,
            I => \N__28912\
        );

    \I__4733\ : Odrv4
    port map (
            O => \N__28912\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__28909\,
            I => \N__28906\
        );

    \I__4731\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28903\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__28903\,
            I => \N__28900\
        );

    \I__4729\ : Odrv12
    port map (
            O => \N__28900\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__4728\ : CascadeMux
    port map (
            O => \N__28897\,
            I => \N__28894\
        );

    \I__4727\ : InMux
    port map (
            O => \N__28894\,
            I => \N__28891\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__28891\,
            I => \N__28888\
        );

    \I__4725\ : Span4Mux_h
    port map (
            O => \N__28888\,
            I => \N__28885\
        );

    \I__4724\ : Odrv4
    port map (
            O => \N__28885\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__28882\,
            I => \N__28879\
        );

    \I__4722\ : InMux
    port map (
            O => \N__28879\,
            I => \N__28876\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__28876\,
            I => \N__28873\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__28873\,
            I => \N__28870\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__28870\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__4718\ : CascadeMux
    port map (
            O => \N__28867\,
            I => \N__28864\
        );

    \I__4717\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28861\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__28861\,
            I => \N__28858\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__28858\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__28855\,
            I => \N__28852\
        );

    \I__4713\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28849\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__28849\,
            I => \N__28846\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__28846\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__4710\ : CascadeMux
    port map (
            O => \N__28843\,
            I => \N__28840\
        );

    \I__4709\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28837\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__28837\,
            I => \N__28834\
        );

    \I__4707\ : Odrv4
    port map (
            O => \N__28834\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__4706\ : InMux
    port map (
            O => \N__28831\,
            I => \N__28825\
        );

    \I__4705\ : InMux
    port map (
            O => \N__28830\,
            I => \N__28818\
        );

    \I__4704\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28818\
        );

    \I__4703\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28818\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__28825\,
            I => \N__28815\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__28818\,
            I => \N__28812\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__28815\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__28812\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__4698\ : InMux
    port map (
            O => \N__28807\,
            I => \N__28803\
        );

    \I__4697\ : InMux
    port map (
            O => \N__28806\,
            I => \N__28800\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__28803\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__28800\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4694\ : InMux
    port map (
            O => \N__28795\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__28792\,
            I => \N__28789\
        );

    \I__4692\ : InMux
    port map (
            O => \N__28789\,
            I => \N__28786\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__28786\,
            I => \N__28783\
        );

    \I__4690\ : Odrv4
    port map (
            O => \N__28783\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19\
        );

    \I__4689\ : CascadeMux
    port map (
            O => \N__28780\,
            I => \N__28777\
        );

    \I__4688\ : InMux
    port map (
            O => \N__28777\,
            I => \N__28774\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__28774\,
            I => \N__28771\
        );

    \I__4686\ : Odrv4
    port map (
            O => \N__28771\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__4685\ : CascadeMux
    port map (
            O => \N__28768\,
            I => \N__28765\
        );

    \I__4684\ : InMux
    port map (
            O => \N__28765\,
            I => \N__28762\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__28762\,
            I => \N__28759\
        );

    \I__4682\ : Span4Mux_h
    port map (
            O => \N__28759\,
            I => \N__28756\
        );

    \I__4681\ : Odrv4
    port map (
            O => \N__28756\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__28753\,
            I => \N__28750\
        );

    \I__4679\ : InMux
    port map (
            O => \N__28750\,
            I => \N__28747\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__28747\,
            I => \N__28744\
        );

    \I__4677\ : Span4Mux_h
    port map (
            O => \N__28744\,
            I => \N__28741\
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__28741\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__28738\,
            I => \N__28735\
        );

    \I__4674\ : InMux
    port map (
            O => \N__28735\,
            I => \N__28732\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__28732\,
            I => \N__28729\
        );

    \I__4672\ : Span4Mux_v
    port map (
            O => \N__28729\,
            I => \N__28726\
        );

    \I__4671\ : Odrv4
    port map (
            O => \N__28726\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__28723\,
            I => \N__28720\
        );

    \I__4669\ : InMux
    port map (
            O => \N__28720\,
            I => \N__28717\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__28717\,
            I => \N__28714\
        );

    \I__4667\ : Odrv4
    port map (
            O => \N__28714\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__28711\,
            I => \N__28708\
        );

    \I__4665\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28705\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28702\
        );

    \I__4663\ : Span4Mux_h
    port map (
            O => \N__28702\,
            I => \N__28699\
        );

    \I__4662\ : Odrv4
    port map (
            O => \N__28699\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__28696\,
            I => \N__28693\
        );

    \I__4660\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28690\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__28690\,
            I => \N__28687\
        );

    \I__4658\ : Odrv12
    port map (
            O => \N__28687\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\
        );

    \I__4657\ : CascadeMux
    port map (
            O => \N__28684\,
            I => \N__28681\
        );

    \I__4656\ : InMux
    port map (
            O => \N__28681\,
            I => \N__28678\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__28678\,
            I => \N__28675\
        );

    \I__4654\ : Span4Mux_h
    port map (
            O => \N__28675\,
            I => \N__28672\
        );

    \I__4653\ : Odrv4
    port map (
            O => \N__28672\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__4652\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28666\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__28666\,
            I => \N__28663\
        );

    \I__4650\ : Span4Mux_h
    port map (
            O => \N__28663\,
            I => \N__28659\
        );

    \I__4649\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28656\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__28659\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__28656\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4646\ : CascadeMux
    port map (
            O => \N__28651\,
            I => \N__28648\
        );

    \I__4645\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28645\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__28645\,
            I => \N__28642\
        );

    \I__4643\ : Span4Mux_h
    port map (
            O => \N__28642\,
            I => \N__28639\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__28639\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11\
        );

    \I__4641\ : InMux
    port map (
            O => \N__28636\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__4640\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28629\
        );

    \I__4639\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28626\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__28629\,
            I => \N__28623\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__28626\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__28623\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4635\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28615\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__28615\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12\
        );

    \I__4633\ : InMux
    port map (
            O => \N__28612\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__4632\ : InMux
    port map (
            O => \N__28609\,
            I => \N__28605\
        );

    \I__4631\ : InMux
    port map (
            O => \N__28608\,
            I => \N__28602\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__28605\,
            I => \N__28599\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__28602\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__28599\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4627\ : CascadeMux
    port map (
            O => \N__28594\,
            I => \N__28591\
        );

    \I__4626\ : InMux
    port map (
            O => \N__28591\,
            I => \N__28588\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__28588\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13\
        );

    \I__4624\ : InMux
    port map (
            O => \N__28585\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__4623\ : InMux
    port map (
            O => \N__28582\,
            I => \N__28578\
        );

    \I__4622\ : InMux
    port map (
            O => \N__28581\,
            I => \N__28575\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__28578\,
            I => \N__28572\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__28575\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__28572\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4618\ : InMux
    port map (
            O => \N__28567\,
            I => \N__28564\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__28564\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14\
        );

    \I__4616\ : InMux
    port map (
            O => \N__28561\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__4615\ : InMux
    port map (
            O => \N__28558\,
            I => \N__28554\
        );

    \I__4614\ : InMux
    port map (
            O => \N__28557\,
            I => \N__28551\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__28554\,
            I => \N__28548\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__28551\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4611\ : Odrv4
    port map (
            O => \N__28548\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__28543\,
            I => \N__28540\
        );

    \I__4609\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28537\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__28537\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15\
        );

    \I__4607\ : InMux
    port map (
            O => \N__28534\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__4606\ : InMux
    port map (
            O => \N__28531\,
            I => \N__28527\
        );

    \I__4605\ : InMux
    port map (
            O => \N__28530\,
            I => \N__28524\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__28527\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__28524\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4602\ : InMux
    port map (
            O => \N__28519\,
            I => \N__28516\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__28516\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16\
        );

    \I__4600\ : InMux
    port map (
            O => \N__28513\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__4599\ : InMux
    port map (
            O => \N__28510\,
            I => \N__28506\
        );

    \I__4598\ : InMux
    port map (
            O => \N__28509\,
            I => \N__28503\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__28506\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__28503\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__28498\,
            I => \N__28495\
        );

    \I__4594\ : InMux
    port map (
            O => \N__28495\,
            I => \N__28492\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__28492\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17\
        );

    \I__4592\ : InMux
    port map (
            O => \N__28489\,
            I => \bfn_11_20_0_\
        );

    \I__4591\ : InMux
    port map (
            O => \N__28486\,
            I => \N__28482\
        );

    \I__4590\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28479\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__28482\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__28479\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4587\ : InMux
    port map (
            O => \N__28474\,
            I => \N__28471\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__28471\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18\
        );

    \I__4585\ : InMux
    port map (
            O => \N__28468\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__28465\,
            I => \N__28462\
        );

    \I__4583\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28458\
        );

    \I__4582\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28455\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__28458\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__28455\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4579\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28447\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__28447\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3\
        );

    \I__4577\ : InMux
    port map (
            O => \N__28444\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__4576\ : InMux
    port map (
            O => \N__28441\,
            I => \N__28437\
        );

    \I__4575\ : InMux
    port map (
            O => \N__28440\,
            I => \N__28434\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__28437\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__28434\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__28429\,
            I => \N__28426\
        );

    \I__4571\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28423\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__28423\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4\
        );

    \I__4569\ : InMux
    port map (
            O => \N__28420\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__4568\ : InMux
    port map (
            O => \N__28417\,
            I => \N__28413\
        );

    \I__4567\ : InMux
    port map (
            O => \N__28416\,
            I => \N__28410\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__28413\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__28410\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__4564\ : InMux
    port map (
            O => \N__28405\,
            I => \N__28402\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__28402\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5\
        );

    \I__4562\ : InMux
    port map (
            O => \N__28399\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__4561\ : InMux
    port map (
            O => \N__28396\,
            I => \N__28392\
        );

    \I__4560\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28389\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__28392\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__28389\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__28384\,
            I => \N__28381\
        );

    \I__4556\ : InMux
    port map (
            O => \N__28381\,
            I => \N__28378\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__28378\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6\
        );

    \I__4554\ : InMux
    port map (
            O => \N__28375\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__4553\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28368\
        );

    \I__4552\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28365\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__28368\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__28365\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__4549\ : InMux
    port map (
            O => \N__28360\,
            I => \N__28357\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__28357\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7\
        );

    \I__4547\ : InMux
    port map (
            O => \N__28354\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__4546\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28347\
        );

    \I__4545\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28344\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__28347\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__28344\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__28339\,
            I => \N__28336\
        );

    \I__4541\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28333\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__28333\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8\
        );

    \I__4539\ : InMux
    port map (
            O => \N__28330\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__4538\ : InMux
    port map (
            O => \N__28327\,
            I => \N__28324\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__28324\,
            I => \N__28320\
        );

    \I__4536\ : InMux
    port map (
            O => \N__28323\,
            I => \N__28317\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__28320\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__28317\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4533\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28309\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__28309\,
            I => \N__28306\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__28306\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9\
        );

    \I__4530\ : InMux
    port map (
            O => \N__28303\,
            I => \bfn_11_19_0_\
        );

    \I__4529\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28297\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28293\
        );

    \I__4527\ : InMux
    port map (
            O => \N__28296\,
            I => \N__28290\
        );

    \I__4526\ : Odrv4
    port map (
            O => \N__28293\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__28290\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4524\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28282\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__28282\,
            I => \N__28279\
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__28279\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10\
        );

    \I__4521\ : InMux
    port map (
            O => \N__28276\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__4520\ : InMux
    port map (
            O => \N__28273\,
            I => \N__28270\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__28270\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__4518\ : CascadeMux
    port map (
            O => \N__28267\,
            I => \N__28264\
        );

    \I__4517\ : InMux
    port map (
            O => \N__28264\,
            I => \N__28261\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__28261\,
            I => \N__28256\
        );

    \I__4515\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28253\
        );

    \I__4514\ : InMux
    port map (
            O => \N__28259\,
            I => \N__28250\
        );

    \I__4513\ : Span4Mux_h
    port map (
            O => \N__28256\,
            I => \N__28247\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__28253\,
            I => \N__28244\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__28250\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__28247\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__28244\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4508\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28233\
        );

    \I__4507\ : InMux
    port map (
            O => \N__28236\,
            I => \N__28230\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__28233\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__28230\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4504\ : CascadeMux
    port map (
            O => \N__28225\,
            I => \N__28222\
        );

    \I__4503\ : InMux
    port map (
            O => \N__28222\,
            I => \N__28219\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__28219\,
            I => \N__28216\
        );

    \I__4501\ : Odrv4
    port map (
            O => \N__28216\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2\
        );

    \I__4500\ : InMux
    port map (
            O => \N__28213\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__4499\ : InMux
    port map (
            O => \N__28210\,
            I => \N__28207\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__28207\,
            I => \N__28204\
        );

    \I__4497\ : Span4Mux_h
    port map (
            O => \N__28204\,
            I => \N__28199\
        );

    \I__4496\ : InMux
    port map (
            O => \N__28203\,
            I => \N__28196\
        );

    \I__4495\ : InMux
    port map (
            O => \N__28202\,
            I => \N__28193\
        );

    \I__4494\ : Odrv4
    port map (
            O => \N__28199\,
            I => measured_delay_tr_12
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__28196\,
            I => measured_delay_tr_12
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__28193\,
            I => measured_delay_tr_12
        );

    \I__4491\ : InMux
    port map (
            O => \N__28186\,
            I => \N__28183\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__28183\,
            I => \N__28180\
        );

    \I__4489\ : Span4Mux_h
    port map (
            O => \N__28180\,
            I => \N__28175\
        );

    \I__4488\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28172\
        );

    \I__4487\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28169\
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__28175\,
            I => measured_delay_tr_11
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__28172\,
            I => measured_delay_tr_11
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__28169\,
            I => measured_delay_tr_11
        );

    \I__4483\ : InMux
    port map (
            O => \N__28162\,
            I => \N__28159\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__28159\,
            I => \N__28155\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__28158\,
            I => \N__28151\
        );

    \I__4480\ : Span4Mux_v
    port map (
            O => \N__28155\,
            I => \N__28148\
        );

    \I__4479\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28145\
        );

    \I__4478\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28142\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__28148\,
            I => measured_delay_tr_13
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__28145\,
            I => measured_delay_tr_13
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__28142\,
            I => measured_delay_tr_13
        );

    \I__4474\ : InMux
    port map (
            O => \N__28135\,
            I => \N__28132\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__28132\,
            I => \N__28128\
        );

    \I__4472\ : InMux
    port map (
            O => \N__28131\,
            I => \N__28124\
        );

    \I__4471\ : Span4Mux_v
    port map (
            O => \N__28128\,
            I => \N__28121\
        );

    \I__4470\ : InMux
    port map (
            O => \N__28127\,
            I => \N__28118\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__28124\,
            I => \N__28115\
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__28121\,
            I => measured_delay_tr_10
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__28118\,
            I => measured_delay_tr_10
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__28115\,
            I => measured_delay_tr_10
        );

    \I__4465\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28105\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__28105\,
            I => \N__28102\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__28102\,
            I => \N__28096\
        );

    \I__4462\ : InMux
    port map (
            O => \N__28101\,
            I => \N__28093\
        );

    \I__4461\ : InMux
    port map (
            O => \N__28100\,
            I => \N__28088\
        );

    \I__4460\ : InMux
    port map (
            O => \N__28099\,
            I => \N__28088\
        );

    \I__4459\ : Odrv4
    port map (
            O => \N__28096\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__28093\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__28088\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__4456\ : InMux
    port map (
            O => \N__28081\,
            I => \N__28077\
        );

    \I__4455\ : InMux
    port map (
            O => \N__28080\,
            I => \N__28074\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__28077\,
            I => \N__28071\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__28074\,
            I => \N__28068\
        );

    \I__4452\ : Span4Mux_h
    port map (
            O => \N__28071\,
            I => \N__28061\
        );

    \I__4451\ : Span4Mux_v
    port map (
            O => \N__28068\,
            I => \N__28061\
        );

    \I__4450\ : InMux
    port map (
            O => \N__28067\,
            I => \N__28058\
        );

    \I__4449\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28055\
        );

    \I__4448\ : Span4Mux_v
    port map (
            O => \N__28061\,
            I => \N__28052\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__28058\,
            I => measured_delay_tr_16
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__28055\,
            I => measured_delay_tr_16
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__28052\,
            I => measured_delay_tr_16
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__28045\,
            I => \N__28042\
        );

    \I__4443\ : InMux
    port map (
            O => \N__28042\,
            I => \N__28039\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__28039\,
            I => \N__28036\
        );

    \I__4441\ : Odrv12
    port map (
            O => \N__28036\,
            I => \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__4440\ : InMux
    port map (
            O => \N__28033\,
            I => \N__28030\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__28030\,
            I => \N__28026\
        );

    \I__4438\ : InMux
    port map (
            O => \N__28029\,
            I => \N__28023\
        );

    \I__4437\ : Span4Mux_h
    port map (
            O => \N__28026\,
            I => \N__28020\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__28023\,
            I => \N__28016\
        );

    \I__4435\ : Span4Mux_v
    port map (
            O => \N__28020\,
            I => \N__28013\
        );

    \I__4434\ : InMux
    port map (
            O => \N__28019\,
            I => \N__28010\
        );

    \I__4433\ : Span4Mux_v
    port map (
            O => \N__28016\,
            I => \N__28007\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__28013\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__28010\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4430\ : Odrv4
    port map (
            O => \N__28007\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__4429\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27996\
        );

    \I__4428\ : InMux
    port map (
            O => \N__27999\,
            I => \N__27993\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__27996\,
            I => \N__27990\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__27993\,
            I => \N__27985\
        );

    \I__4425\ : Span4Mux_v
    port map (
            O => \N__27990\,
            I => \N__27982\
        );

    \I__4424\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27979\
        );

    \I__4423\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27976\
        );

    \I__4422\ : Span4Mux_h
    port map (
            O => \N__27985\,
            I => \N__27971\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__27982\,
            I => \N__27971\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__27979\,
            I => \N__27968\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__27976\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__27971\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__4417\ : Odrv12
    port map (
            O => \N__27968\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__4416\ : InMux
    port map (
            O => \N__27961\,
            I => \N__27958\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__27958\,
            I => \N__27955\
        );

    \I__4414\ : Span4Mux_h
    port map (
            O => \N__27955\,
            I => \N__27952\
        );

    \I__4413\ : Odrv4
    port map (
            O => \N__27952\,
            I => \phase_controller_inst2.start_timer_hc_RNO_0_0\
        );

    \I__4412\ : InMux
    port map (
            O => \N__27949\,
            I => \N__27945\
        );

    \I__4411\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27942\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__27945\,
            I => \N__27938\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__27942\,
            I => \N__27935\
        );

    \I__4408\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27932\
        );

    \I__4407\ : Span12Mux_v
    port map (
            O => \N__27938\,
            I => \N__27929\
        );

    \I__4406\ : Span4Mux_v
    port map (
            O => \N__27935\,
            I => \N__27926\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__27932\,
            I => measured_delay_tr_4
        );

    \I__4404\ : Odrv12
    port map (
            O => \N__27929\,
            I => measured_delay_tr_4
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__27926\,
            I => measured_delay_tr_4
        );

    \I__4402\ : CascadeMux
    port map (
            O => \N__27919\,
            I => \N__27916\
        );

    \I__4401\ : InMux
    port map (
            O => \N__27916\,
            I => \N__27912\
        );

    \I__4400\ : InMux
    port map (
            O => \N__27915\,
            I => \N__27909\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__27912\,
            I => \N__27905\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__27909\,
            I => \N__27902\
        );

    \I__4397\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27899\
        );

    \I__4396\ : Span4Mux_v
    port map (
            O => \N__27905\,
            I => \N__27896\
        );

    \I__4395\ : Span4Mux_v
    port map (
            O => \N__27902\,
            I => \N__27893\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__27899\,
            I => measured_delay_tr_9
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__27896\,
            I => measured_delay_tr_9
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__27893\,
            I => measured_delay_tr_9
        );

    \I__4391\ : CascadeMux
    port map (
            O => \N__27886\,
            I => \N__27883\
        );

    \I__4390\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27878\
        );

    \I__4389\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27875\
        );

    \I__4388\ : CascadeMux
    port map (
            O => \N__27881\,
            I => \N__27872\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__27878\,
            I => \N__27867\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__27875\,
            I => \N__27867\
        );

    \I__4385\ : InMux
    port map (
            O => \N__27872\,
            I => \N__27864\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__27867\,
            I => \N__27861\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__27864\,
            I => measured_delay_tr_3
        );

    \I__4382\ : Odrv4
    port map (
            O => \N__27861\,
            I => measured_delay_tr_3
        );

    \I__4381\ : CascadeMux
    port map (
            O => \N__27856\,
            I => \N__27853\
        );

    \I__4380\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27850\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__27850\,
            I => \N__27845\
        );

    \I__4378\ : InMux
    port map (
            O => \N__27849\,
            I => \N__27842\
        );

    \I__4377\ : InMux
    port map (
            O => \N__27848\,
            I => \N__27839\
        );

    \I__4376\ : Span4Mux_h
    port map (
            O => \N__27845\,
            I => \N__27834\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__27842\,
            I => \N__27834\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__27839\,
            I => measured_delay_tr_2
        );

    \I__4373\ : Odrv4
    port map (
            O => \N__27834\,
            I => measured_delay_tr_2
        );

    \I__4372\ : InMux
    port map (
            O => \N__27829\,
            I => \N__27825\
        );

    \I__4371\ : InMux
    port map (
            O => \N__27828\,
            I => \N__27822\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__27825\,
            I => \N__27818\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__27822\,
            I => \N__27815\
        );

    \I__4368\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27812\
        );

    \I__4367\ : Span4Mux_v
    port map (
            O => \N__27818\,
            I => \N__27809\
        );

    \I__4366\ : Span4Mux_h
    port map (
            O => \N__27815\,
            I => \N__27804\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__27812\,
            I => \N__27804\
        );

    \I__4364\ : Odrv4
    port map (
            O => \N__27809\,
            I => measured_delay_tr_6
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__27804\,
            I => measured_delay_tr_6
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__27799\,
            I => \N__27796\
        );

    \I__4361\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27793\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__27793\,
            I => \N__27789\
        );

    \I__4359\ : CascadeMux
    port map (
            O => \N__27792\,
            I => \N__27786\
        );

    \I__4358\ : Span4Mux_h
    port map (
            O => \N__27789\,
            I => \N__27783\
        );

    \I__4357\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27780\
        );

    \I__4356\ : Odrv4
    port map (
            O => \N__27783\,
            I => measured_delay_tr_1
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__27780\,
            I => measured_delay_tr_1
        );

    \I__4354\ : InMux
    port map (
            O => \N__27775\,
            I => \N__27772\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__27772\,
            I => \N__27767\
        );

    \I__4352\ : InMux
    port map (
            O => \N__27771\,
            I => \N__27760\
        );

    \I__4351\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27760\
        );

    \I__4350\ : Span4Mux_v
    port map (
            O => \N__27767\,
            I => \N__27757\
        );

    \I__4349\ : InMux
    port map (
            O => \N__27766\,
            I => \N__27752\
        );

    \I__4348\ : InMux
    port map (
            O => \N__27765\,
            I => \N__27752\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__27760\,
            I => \N__27749\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__27757\,
            I => measured_delay_tr_14
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__27752\,
            I => measured_delay_tr_14
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__27749\,
            I => measured_delay_tr_14
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__27742\,
            I => \N__27739\
        );

    \I__4342\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27736\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__27736\,
            I => \N__27733\
        );

    \I__4340\ : Odrv4
    port map (
            O => \N__27733\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__27730\,
            I => \N__27727\
        );

    \I__4338\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27724\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__27724\,
            I => \N__27721\
        );

    \I__4336\ : Span4Mux_v
    port map (
            O => \N__27721\,
            I => \N__27718\
        );

    \I__4335\ : Odrv4
    port map (
            O => \N__27718\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__4334\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27712\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__27712\,
            I => \N__27707\
        );

    \I__4332\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27703\
        );

    \I__4331\ : CascadeMux
    port map (
            O => \N__27710\,
            I => \N__27700\
        );

    \I__4330\ : Span4Mux_h
    port map (
            O => \N__27707\,
            I => \N__27697\
        );

    \I__4329\ : InMux
    port map (
            O => \N__27706\,
            I => \N__27694\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__27703\,
            I => \N__27691\
        );

    \I__4327\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27688\
        );

    \I__4326\ : Span4Mux_v
    port map (
            O => \N__27697\,
            I => \N__27685\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__27694\,
            I => \N__27680\
        );

    \I__4324\ : Span4Mux_v
    port map (
            O => \N__27691\,
            I => \N__27680\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__27688\,
            I => measured_delay_tr_8
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__27685\,
            I => measured_delay_tr_8
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__27680\,
            I => measured_delay_tr_8
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__27673\,
            I => \N__27670\
        );

    \I__4319\ : InMux
    port map (
            O => \N__27670\,
            I => \N__27667\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__27667\,
            I => \N__27664\
        );

    \I__4317\ : Span4Mux_h
    port map (
            O => \N__27664\,
            I => \N__27661\
        );

    \I__4316\ : Odrv4
    port map (
            O => \N__27661\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__4315\ : CascadeMux
    port map (
            O => \N__27658\,
            I => \N__27655\
        );

    \I__4314\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27652\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__27652\,
            I => \N__27649\
        );

    \I__4312\ : Odrv4
    port map (
            O => \N__27649\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__4311\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27643\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__27643\,
            I => \N__27639\
        );

    \I__4309\ : InMux
    port map (
            O => \N__27642\,
            I => \N__27636\
        );

    \I__4308\ : Span4Mux_v
    port map (
            O => \N__27639\,
            I => \N__27630\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__27636\,
            I => \N__27630\
        );

    \I__4306\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27627\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__27630\,
            I => \N__27624\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__27627\,
            I => measured_delay_tr_5
        );

    \I__4303\ : Odrv4
    port map (
            O => \N__27624\,
            I => measured_delay_tr_5
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__27619\,
            I => \N__27616\
        );

    \I__4301\ : InMux
    port map (
            O => \N__27616\,
            I => \N__27613\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__27613\,
            I => \N__27610\
        );

    \I__4299\ : Span4Mux_h
    port map (
            O => \N__27610\,
            I => \N__27607\
        );

    \I__4298\ : Odrv4
    port map (
            O => \N__27607\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__4297\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27601\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__27601\,
            I => \N__27598\
        );

    \I__4295\ : Odrv12
    port map (
            O => \N__27598\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__27595\,
            I => \N__27592\
        );

    \I__4293\ : InMux
    port map (
            O => \N__27592\,
            I => \N__27589\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__27589\,
            I => \N__27586\
        );

    \I__4291\ : Odrv12
    port map (
            O => \N__27586\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__27583\,
            I => \N__27580\
        );

    \I__4289\ : InMux
    port map (
            O => \N__27580\,
            I => \N__27577\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__27577\,
            I => \N__27574\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__27574\,
            I => \N__27571\
        );

    \I__4286\ : Odrv4
    port map (
            O => \N__27571\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__4285\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27563\
        );

    \I__4284\ : CascadeMux
    port map (
            O => \N__27567\,
            I => \N__27559\
        );

    \I__4283\ : InMux
    port map (
            O => \N__27566\,
            I => \N__27556\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__27563\,
            I => \N__27553\
        );

    \I__4281\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27550\
        );

    \I__4280\ : InMux
    port map (
            O => \N__27559\,
            I => \N__27547\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__27556\,
            I => \N__27542\
        );

    \I__4278\ : Span4Mux_v
    port map (
            O => \N__27553\,
            I => \N__27542\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__27550\,
            I => \N__27539\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__27547\,
            I => \N__27534\
        );

    \I__4275\ : Span4Mux_v
    port map (
            O => \N__27542\,
            I => \N__27534\
        );

    \I__4274\ : Span4Mux_v
    port map (
            O => \N__27539\,
            I => \N__27531\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__27534\,
            I => measured_delay_tr_7
        );

    \I__4272\ : Odrv4
    port map (
            O => \N__27531\,
            I => measured_delay_tr_7
        );

    \I__4271\ : CascadeMux
    port map (
            O => \N__27526\,
            I => \N__27523\
        );

    \I__4270\ : InMux
    port map (
            O => \N__27523\,
            I => \N__27520\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__27520\,
            I => \N__27517\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__27517\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__4267\ : CascadeMux
    port map (
            O => \N__27514\,
            I => \N__27511\
        );

    \I__4266\ : InMux
    port map (
            O => \N__27511\,
            I => \N__27508\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__27508\,
            I => \N__27505\
        );

    \I__4264\ : Odrv4
    port map (
            O => \N__27505\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__4263\ : InMux
    port map (
            O => \N__27502\,
            I => \N__27498\
        );

    \I__4262\ : InMux
    port map (
            O => \N__27501\,
            I => \N__27495\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__27498\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__27495\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4259\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27487\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__27487\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\
        );

    \I__4257\ : InMux
    port map (
            O => \N__27484\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__4256\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27477\
        );

    \I__4255\ : InMux
    port map (
            O => \N__27480\,
            I => \N__27474\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__27477\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__27474\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4252\ : InMux
    port map (
            O => \N__27469\,
            I => \N__27466\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__27466\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\
        );

    \I__4250\ : InMux
    port map (
            O => \N__27463\,
            I => \bfn_10_26_0_\
        );

    \I__4249\ : InMux
    port map (
            O => \N__27460\,
            I => \N__27456\
        );

    \I__4248\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27453\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__27456\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__27453\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4245\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27445\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__27445\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\
        );

    \I__4243\ : InMux
    port map (
            O => \N__27442\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__4242\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27435\
        );

    \I__4241\ : InMux
    port map (
            O => \N__27438\,
            I => \N__27432\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__27435\,
            I => \N__27429\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__27432\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4238\ : Odrv4
    port map (
            O => \N__27429\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4237\ : InMux
    port map (
            O => \N__27424\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__4236\ : InMux
    port map (
            O => \N__27421\,
            I => \N__27418\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__27418\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\
        );

    \I__4234\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27412\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__27412\,
            I => \N__27409\
        );

    \I__4232\ : Span12Mux_h
    port map (
            O => \N__27409\,
            I => \N__27406\
        );

    \I__4231\ : Odrv12
    port map (
            O => \N__27406\,
            I => delay_hc_input_c
        );

    \I__4230\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27400\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__27400\,
            I => delay_hc_d1
        );

    \I__4228\ : InMux
    port map (
            O => \N__27397\,
            I => \N__27394\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__27394\,
            I => \N__27389\
        );

    \I__4226\ : InMux
    port map (
            O => \N__27393\,
            I => \N__27386\
        );

    \I__4225\ : InMux
    port map (
            O => \N__27392\,
            I => \N__27382\
        );

    \I__4224\ : Span4Mux_h
    port map (
            O => \N__27389\,
            I => \N__27379\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__27386\,
            I => \N__27376\
        );

    \I__4222\ : InMux
    port map (
            O => \N__27385\,
            I => \N__27373\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__27382\,
            I => delay_hc_d2
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__27379\,
            I => delay_hc_d2
        );

    \I__4219\ : Odrv4
    port map (
            O => \N__27376\,
            I => delay_hc_d2
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__27373\,
            I => delay_hc_d2
        );

    \I__4217\ : InMux
    port map (
            O => \N__27364\,
            I => \N__27360\
        );

    \I__4216\ : InMux
    port map (
            O => \N__27363\,
            I => \N__27356\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__27360\,
            I => \N__27353\
        );

    \I__4214\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27350\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__27356\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__27353\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__27350\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__4210\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27339\
        );

    \I__4209\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27336\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__27339\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__27336\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__4206\ : InMux
    port map (
            O => \N__27331\,
            I => \N__27328\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__27328\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\
        );

    \I__4204\ : InMux
    port map (
            O => \N__27325\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__4203\ : InMux
    port map (
            O => \N__27322\,
            I => \N__27319\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__27319\,
            I => \N__27315\
        );

    \I__4201\ : InMux
    port map (
            O => \N__27318\,
            I => \N__27312\
        );

    \I__4200\ : Odrv12
    port map (
            O => \N__27315\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__27312\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4198\ : InMux
    port map (
            O => \N__27307\,
            I => \N__27304\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__27304\,
            I => \N__27301\
        );

    \I__4196\ : Odrv4
    port map (
            O => \N__27301\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\
        );

    \I__4195\ : InMux
    port map (
            O => \N__27298\,
            I => \bfn_10_25_0_\
        );

    \I__4194\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27292\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__27292\,
            I => \N__27288\
        );

    \I__4192\ : InMux
    port map (
            O => \N__27291\,
            I => \N__27285\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__27288\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__27285\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4189\ : InMux
    port map (
            O => \N__27280\,
            I => \N__27277\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__27277\,
            I => \N__27274\
        );

    \I__4187\ : Odrv4
    port map (
            O => \N__27274\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\
        );

    \I__4186\ : InMux
    port map (
            O => \N__27271\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__4185\ : InMux
    port map (
            O => \N__27268\,
            I => \N__27264\
        );

    \I__4184\ : InMux
    port map (
            O => \N__27267\,
            I => \N__27261\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__27264\,
            I => \N__27258\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__27261\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4181\ : Odrv4
    port map (
            O => \N__27258\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4180\ : InMux
    port map (
            O => \N__27253\,
            I => \N__27250\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__27250\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\
        );

    \I__4178\ : InMux
    port map (
            O => \N__27247\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__4177\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27240\
        );

    \I__4176\ : InMux
    port map (
            O => \N__27243\,
            I => \N__27237\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__27240\,
            I => \N__27234\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__27237\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__27234\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4172\ : InMux
    port map (
            O => \N__27229\,
            I => \N__27226\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__27226\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\
        );

    \I__4170\ : InMux
    port map (
            O => \N__27223\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__4169\ : InMux
    port map (
            O => \N__27220\,
            I => \N__27216\
        );

    \I__4168\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27213\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__27216\,
            I => \N__27210\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__27213\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__27210\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4164\ : InMux
    port map (
            O => \N__27205\,
            I => \N__27202\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__27202\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\
        );

    \I__4162\ : InMux
    port map (
            O => \N__27199\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__4161\ : InMux
    port map (
            O => \N__27196\,
            I => \N__27192\
        );

    \I__4160\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27189\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__27192\,
            I => \N__27186\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__27189\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4157\ : Odrv4
    port map (
            O => \N__27186\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4156\ : InMux
    port map (
            O => \N__27181\,
            I => \N__27178\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__27178\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\
        );

    \I__4154\ : InMux
    port map (
            O => \N__27175\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__4153\ : InMux
    port map (
            O => \N__27172\,
            I => \N__27168\
        );

    \I__4152\ : InMux
    port map (
            O => \N__27171\,
            I => \N__27165\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__27168\,
            I => \N__27162\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__27165\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__27162\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4148\ : InMux
    port map (
            O => \N__27157\,
            I => \N__27154\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__27154\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\
        );

    \I__4146\ : InMux
    port map (
            O => \N__27151\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__4145\ : InMux
    port map (
            O => \N__27148\,
            I => \N__27145\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__27145\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__27142\,
            I => \N__27138\
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__27141\,
            I => \N__27135\
        );

    \I__4141\ : InMux
    port map (
            O => \N__27138\,
            I => \N__27132\
        );

    \I__4140\ : InMux
    port map (
            O => \N__27135\,
            I => \N__27129\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__27132\,
            I => \N__27123\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__27129\,
            I => \N__27123\
        );

    \I__4137\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27120\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__27123\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__27120\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4134\ : InMux
    port map (
            O => \N__27115\,
            I => \N__27111\
        );

    \I__4133\ : InMux
    port map (
            O => \N__27114\,
            I => \N__27108\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__27111\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__27108\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4130\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27100\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__27100\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\
        );

    \I__4128\ : InMux
    port map (
            O => \N__27097\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__4127\ : InMux
    port map (
            O => \N__27094\,
            I => \N__27091\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__27091\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\
        );

    \I__4125\ : CascadeMux
    port map (
            O => \N__27088\,
            I => \N__27085\
        );

    \I__4124\ : InMux
    port map (
            O => \N__27085\,
            I => \N__27081\
        );

    \I__4123\ : InMux
    port map (
            O => \N__27084\,
            I => \N__27078\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__27081\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__27078\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4120\ : InMux
    port map (
            O => \N__27073\,
            I => \N__27070\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__27070\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\
        );

    \I__4118\ : InMux
    port map (
            O => \N__27067\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__4117\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27060\
        );

    \I__4116\ : InMux
    port map (
            O => \N__27063\,
            I => \N__27057\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__27060\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__27057\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4113\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27049\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__27049\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\
        );

    \I__4111\ : InMux
    port map (
            O => \N__27046\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__4110\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27039\
        );

    \I__4109\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27036\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__27039\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__27036\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__4106\ : InMux
    port map (
            O => \N__27031\,
            I => \N__27028\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__27028\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\
        );

    \I__4104\ : InMux
    port map (
            O => \N__27025\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__4103\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27018\
        );

    \I__4102\ : InMux
    port map (
            O => \N__27021\,
            I => \N__27015\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__27018\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__27015\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__4099\ : InMux
    port map (
            O => \N__27010\,
            I => \N__27007\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__27007\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\
        );

    \I__4097\ : InMux
    port map (
            O => \N__27004\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__4096\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26997\
        );

    \I__4095\ : InMux
    port map (
            O => \N__27000\,
            I => \N__26994\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__26997\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__26994\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__4092\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26986\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__26986\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26983\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__26980\,
            I => \N__26977\
        );

    \I__4088\ : InMux
    port map (
            O => \N__26977\,
            I => \N__26974\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__26974\,
            I => \N__26971\
        );

    \I__4086\ : Odrv12
    port map (
            O => \N__26971\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26968\,
            I => \N__26965\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__26965\,
            I => \N__26962\
        );

    \I__4083\ : Span4Mux_h
    port map (
            O => \N__26962\,
            I => \N__26959\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__26959\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__26956\,
            I => \N__26953\
        );

    \I__4080\ : InMux
    port map (
            O => \N__26953\,
            I => \N__26950\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__26950\,
            I => \N__26947\
        );

    \I__4078\ : Span4Mux_h
    port map (
            O => \N__26947\,
            I => \N__26944\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__26944\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ1Z_6\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__26941\,
            I => \N__26938\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26935\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__26935\,
            I => \N__26932\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__26932\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__4072\ : InMux
    port map (
            O => \N__26929\,
            I => \N__26926\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__26926\,
            I => \N__26923\
        );

    \I__4070\ : Span4Mux_h
    port map (
            O => \N__26923\,
            I => \N__26920\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__26920\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_0\
        );

    \I__4068\ : CascadeMux
    port map (
            O => \N__26917\,
            I => \N__26914\
        );

    \I__4067\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26911\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__26911\,
            I => \N__26908\
        );

    \I__4065\ : Odrv12
    port map (
            O => \N__26908\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__26905\,
            I => \N__26902\
        );

    \I__4063\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26899\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__26899\,
            I => \N__26896\
        );

    \I__4061\ : Span4Mux_h
    port map (
            O => \N__26896\,
            I => \N__26893\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__26893\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__26890\,
            I => \N__26887\
        );

    \I__4058\ : InMux
    port map (
            O => \N__26887\,
            I => \N__26884\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__26884\,
            I => \N__26881\
        );

    \I__4056\ : Span4Mux_v
    port map (
            O => \N__26881\,
            I => \N__26878\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__26878\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26875\,
            I => \N__26872\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26872\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\
        );

    \I__4052\ : InMux
    port map (
            O => \N__26869\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__4051\ : InMux
    port map (
            O => \N__26866\,
            I => \N__26863\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__26863\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__4049\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26857\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__26857\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__4047\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26851\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__26851\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__4045\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26845\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__26845\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__4043\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26839\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__26839\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__4041\ : InMux
    port map (
            O => \N__26836\,
            I => \N__26833\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__26833\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__4039\ : InMux
    port map (
            O => \N__26830\,
            I => \N__26827\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__26827\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\
        );

    \I__4037\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26821\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__26821\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\
        );

    \I__4035\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26815\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__26815\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\
        );

    \I__4033\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26809\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__26809\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__4031\ : InMux
    port map (
            O => \N__26806\,
            I => \N__26803\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__26803\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__4029\ : InMux
    port map (
            O => \N__26800\,
            I => \N__26797\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__26797\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__4027\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26791\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__26791\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__4025\ : InMux
    port map (
            O => \N__26788\,
            I => \N__26785\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__26785\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__4023\ : InMux
    port map (
            O => \N__26782\,
            I => \N__26779\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__26779\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__4021\ : InMux
    port map (
            O => \N__26776\,
            I => \N__26773\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__26773\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__4019\ : InMux
    port map (
            O => \N__26770\,
            I => \N__26767\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__26767\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__26764\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_\
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__26761\,
            I => \N__26756\
        );

    \I__4015\ : CascadeMux
    port map (
            O => \N__26760\,
            I => \N__26751\
        );

    \I__4014\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26746\
        );

    \I__4013\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26733\
        );

    \I__4012\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26733\
        );

    \I__4011\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26733\
        );

    \I__4010\ : InMux
    port map (
            O => \N__26751\,
            I => \N__26733\
        );

    \I__4009\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26733\
        );

    \I__4008\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26733\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26725\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__26733\,
            I => \N__26722\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26719\
        );

    \I__4004\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26706\
        );

    \I__4003\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26706\
        );

    \I__4002\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26706\
        );

    \I__4001\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26706\
        );

    \I__4000\ : Span4Mux_v
    port map (
            O => \N__26725\,
            I => \N__26699\
        );

    \I__3999\ : Span4Mux_h
    port map (
            O => \N__26722\,
            I => \N__26699\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__26719\,
            I => \N__26699\
        );

    \I__3997\ : InMux
    port map (
            O => \N__26718\,
            I => \N__26690\
        );

    \I__3996\ : InMux
    port map (
            O => \N__26717\,
            I => \N__26690\
        );

    \I__3995\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26690\
        );

    \I__3994\ : InMux
    port map (
            O => \N__26715\,
            I => \N__26690\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__26706\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__26699\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__26690\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__26683\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\
        );

    \I__3989\ : InMux
    port map (
            O => \N__26680\,
            I => \N__26677\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__26677\,
            I => \N__26667\
        );

    \I__3987\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26658\
        );

    \I__3986\ : InMux
    port map (
            O => \N__26675\,
            I => \N__26658\
        );

    \I__3985\ : InMux
    port map (
            O => \N__26674\,
            I => \N__26658\
        );

    \I__3984\ : InMux
    port map (
            O => \N__26673\,
            I => \N__26658\
        );

    \I__3983\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26655\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__26671\,
            I => \N__26652\
        );

    \I__3981\ : CascadeMux
    port map (
            O => \N__26670\,
            I => \N__26649\
        );

    \I__3980\ : Span4Mux_h
    port map (
            O => \N__26667\,
            I => \N__26641\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__26658\,
            I => \N__26641\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__26655\,
            I => \N__26641\
        );

    \I__3977\ : InMux
    port map (
            O => \N__26652\,
            I => \N__26631\
        );

    \I__3976\ : InMux
    port map (
            O => \N__26649\,
            I => \N__26631\
        );

    \I__3975\ : InMux
    port map (
            O => \N__26648\,
            I => \N__26631\
        );

    \I__3974\ : Span4Mux_v
    port map (
            O => \N__26641\,
            I => \N__26628\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26640\,
            I => \N__26621\
        );

    \I__3972\ : InMux
    port map (
            O => \N__26639\,
            I => \N__26621\
        );

    \I__3971\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26621\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__26631\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__26628\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__26621\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__3967\ : InMux
    port map (
            O => \N__26614\,
            I => \N__26611\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__26611\,
            I => \N__26608\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__26608\,
            I => \N__26605\
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__26605\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\
        );

    \I__3963\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26599\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__26599\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__26596\,
            I => \N__26593\
        );

    \I__3960\ : InMux
    port map (
            O => \N__26593\,
            I => \N__26590\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__26590\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\
        );

    \I__3958\ : InMux
    port map (
            O => \N__26587\,
            I => \N__26584\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__26584\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\
        );

    \I__3956\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26578\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__26578\,
            I => \N__26574\
        );

    \I__3954\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26571\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__26574\,
            I => \phase_controller_inst1.stoper_tr.N_248\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__26571\,
            I => \phase_controller_inst1.stoper_tr.N_248\
        );

    \I__3951\ : CascadeMux
    port map (
            O => \N__26566\,
            I => \phase_controller_inst1.stoper_tr.N_248_cascade_\
        );

    \I__3950\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26557\
        );

    \I__3949\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26557\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__26557\,
            I => \N__26552\
        );

    \I__3947\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26547\
        );

    \I__3946\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26547\
        );

    \I__3945\ : Odrv12
    port map (
            O => \N__26552\,
            I => \phase_controller_inst1.stoper_tr.N_55\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__26547\,
            I => \phase_controller_inst1.stoper_tr.N_55\
        );

    \I__3943\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26539\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__26539\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__3941\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26533\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__26533\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__3939\ : CascadeMux
    port map (
            O => \N__26530\,
            I => \N__26527\
        );

    \I__3938\ : InMux
    port map (
            O => \N__26527\,
            I => \N__26524\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__26524\,
            I => \N__26521\
        );

    \I__3936\ : Odrv4
    port map (
            O => \N__26521\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__26518\,
            I => \N__26515\
        );

    \I__3934\ : InMux
    port map (
            O => \N__26515\,
            I => \N__26512\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__26512\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__3932\ : CascadeMux
    port map (
            O => \N__26509\,
            I => \N__26506\
        );

    \I__3931\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26503\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__26503\,
            I => \N__26500\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__26500\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__26497\,
            I => \N__26494\
        );

    \I__3927\ : InMux
    port map (
            O => \N__26494\,
            I => \N__26491\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__26491\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__26488\,
            I => \N__26485\
        );

    \I__3924\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26482\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__26482\,
            I => \N__26479\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__26479\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__26476\,
            I => \N__26473\
        );

    \I__3920\ : InMux
    port map (
            O => \N__26473\,
            I => \N__26470\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__26470\,
            I => \N__26467\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__26467\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__3917\ : InMux
    port map (
            O => \N__26464\,
            I => \N__26461\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__26461\,
            I => \N__26454\
        );

    \I__3915\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26447\
        );

    \I__3914\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26447\
        );

    \I__3913\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26447\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__26457\,
            I => \N__26443\
        );

    \I__3911\ : Span4Mux_h
    port map (
            O => \N__26454\,
            I => \N__26436\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__26447\,
            I => \N__26433\
        );

    \I__3909\ : InMux
    port map (
            O => \N__26446\,
            I => \N__26430\
        );

    \I__3908\ : InMux
    port map (
            O => \N__26443\,
            I => \N__26419\
        );

    \I__3907\ : InMux
    port map (
            O => \N__26442\,
            I => \N__26419\
        );

    \I__3906\ : InMux
    port map (
            O => \N__26441\,
            I => \N__26419\
        );

    \I__3905\ : InMux
    port map (
            O => \N__26440\,
            I => \N__26419\
        );

    \I__3904\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26419\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__26436\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__26433\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__26430\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__26419\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__3899\ : CascadeMux
    port map (
            O => \N__26410\,
            I => \N__26407\
        );

    \I__3898\ : InMux
    port map (
            O => \N__26407\,
            I => \N__26404\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__26404\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__3896\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26397\
        );

    \I__3895\ : InMux
    port map (
            O => \N__26400\,
            I => \N__26394\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__26397\,
            I => \N__26389\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__26394\,
            I => \N__26389\
        );

    \I__3892\ : Odrv12
    port map (
            O => \N__26389\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__3891\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26381\
        );

    \I__3890\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26378\
        );

    \I__3889\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26375\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__26381\,
            I => \N__26372\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__26378\,
            I => \N__26367\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__26375\,
            I => \N__26367\
        );

    \I__3885\ : Span4Mux_h
    port map (
            O => \N__26372\,
            I => \N__26364\
        );

    \I__3884\ : Span4Mux_v
    port map (
            O => \N__26367\,
            I => \N__26361\
        );

    \I__3883\ : Span4Mux_v
    port map (
            O => \N__26364\,
            I => \N__26358\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__26361\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__26358\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__26353\,
            I => \N__26350\
        );

    \I__3879\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26347\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__26347\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__26344\,
            I => \N__26341\
        );

    \I__3876\ : InMux
    port map (
            O => \N__26341\,
            I => \N__26338\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__26338\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__3874\ : CascadeMux
    port map (
            O => \N__26335\,
            I => \N__26332\
        );

    \I__3873\ : InMux
    port map (
            O => \N__26332\,
            I => \N__26329\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__26329\,
            I => \N__26326\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__26326\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__26323\,
            I => \N__26320\
        );

    \I__3869\ : InMux
    port map (
            O => \N__26320\,
            I => \N__26317\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__26317\,
            I => \N__26314\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__26314\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__26311\,
            I => \N__26308\
        );

    \I__3865\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26305\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__26305\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__26302\,
            I => \N__26299\
        );

    \I__3862\ : InMux
    port map (
            O => \N__26299\,
            I => \N__26296\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__26296\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__3860\ : CascadeMux
    port map (
            O => \N__26293\,
            I => \N__26290\
        );

    \I__3859\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26287\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__26287\,
            I => \N__26284\
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__26284\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__26281\,
            I => \N__26278\
        );

    \I__3855\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26275\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__26275\,
            I => \N__26272\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__26272\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__26269\,
            I => \N__26266\
        );

    \I__3851\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26263\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__26263\,
            I => \N__26260\
        );

    \I__3849\ : Odrv4
    port map (
            O => \N__26260\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__3848\ : CascadeMux
    port map (
            O => \N__26257\,
            I => \N__26254\
        );

    \I__3847\ : InMux
    port map (
            O => \N__26254\,
            I => \N__26251\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__26251\,
            I => \N__26248\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__26248\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__26245\,
            I => \N__26242\
        );

    \I__3843\ : InMux
    port map (
            O => \N__26242\,
            I => \N__26239\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__26239\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__26236\,
            I => \N__26233\
        );

    \I__3840\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26230\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__26230\,
            I => \N__26227\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__26227\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__3837\ : InMux
    port map (
            O => \N__26224\,
            I => \N__26221\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__26221\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__3835\ : CascadeMux
    port map (
            O => \N__26218\,
            I => \N__26212\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__26217\,
            I => \N__26208\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__26216\,
            I => \N__26204\
        );

    \I__3832\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26191\
        );

    \I__3831\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26191\
        );

    \I__3830\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26191\
        );

    \I__3829\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26191\
        );

    \I__3828\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26191\
        );

    \I__3827\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26191\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__26191\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__26188\,
            I => \N__26185\
        );

    \I__3824\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26182\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__26182\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__3822\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26174\
        );

    \I__3821\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26171\
        );

    \I__3820\ : InMux
    port map (
            O => \N__26177\,
            I => \N__26168\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__26174\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__26171\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__26168\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__26161\,
            I => \N__26158\
        );

    \I__3815\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26155\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__26155\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__3813\ : InMux
    port map (
            O => \N__26152\,
            I => \N__26149\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__26149\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__26146\,
            I => \N__26143\
        );

    \I__3810\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26140\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__26140\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__26137\,
            I => \N__26134\
        );

    \I__3807\ : InMux
    port map (
            O => \N__26134\,
            I => \N__26131\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__26131\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__3805\ : InMux
    port map (
            O => \N__26128\,
            I => \N__26125\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__26125\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__3803\ : InMux
    port map (
            O => \N__26122\,
            I => \N__26119\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__26119\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__26116\,
            I => \N__26113\
        );

    \I__3800\ : InMux
    port map (
            O => \N__26113\,
            I => \N__26110\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__26110\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__3798\ : InMux
    port map (
            O => \N__26107\,
            I => \N__26104\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__26104\,
            I => \N__26100\
        );

    \I__3796\ : CascadeMux
    port map (
            O => \N__26103\,
            I => \N__26097\
        );

    \I__3795\ : Span4Mux_v
    port map (
            O => \N__26100\,
            I => \N__26092\
        );

    \I__3794\ : InMux
    port map (
            O => \N__26097\,
            I => \N__26087\
        );

    \I__3793\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26087\
        );

    \I__3792\ : InMux
    port map (
            O => \N__26095\,
            I => \N__26084\
        );

    \I__3791\ : Span4Mux_v
    port map (
            O => \N__26092\,
            I => \N__26079\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__26087\,
            I => \N__26079\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__26084\,
            I => \N__26074\
        );

    \I__3788\ : Span4Mux_v
    port map (
            O => \N__26079\,
            I => \N__26074\
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__26074\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__3786\ : IoInMux
    port map (
            O => \N__26071\,
            I => \N__26068\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__26068\,
            I => \N__26065\
        );

    \I__3784\ : Odrv12
    port map (
            O => \N__26065\,
            I => s3_phy_c
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__26062\,
            I => \N__26058\
        );

    \I__3782\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26055\
        );

    \I__3781\ : InMux
    port map (
            O => \N__26058\,
            I => \N__26052\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__26055\,
            I => \N__26048\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__26052\,
            I => \N__26045\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__26051\,
            I => \N__26042\
        );

    \I__3777\ : Span12Mux_v
    port map (
            O => \N__26048\,
            I => \N__26038\
        );

    \I__3776\ : Span4Mux_v
    port map (
            O => \N__26045\,
            I => \N__26035\
        );

    \I__3775\ : InMux
    port map (
            O => \N__26042\,
            I => \N__26032\
        );

    \I__3774\ : InMux
    port map (
            O => \N__26041\,
            I => \N__26029\
        );

    \I__3773\ : Odrv12
    port map (
            O => \N__26038\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__26035\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__26032\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__26029\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__3769\ : IoInMux
    port map (
            O => \N__26020\,
            I => \N__26017\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__26017\,
            I => \N__26014\
        );

    \I__3767\ : Span4Mux_s1_v
    port map (
            O => \N__26014\,
            I => \N__26011\
        );

    \I__3766\ : Span4Mux_h
    port map (
            O => \N__26011\,
            I => \N__26008\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__26008\,
            I => s2_phy_c
        );

    \I__3764\ : InMux
    port map (
            O => \N__26005\,
            I => \N__26002\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__26002\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__3762\ : InMux
    port map (
            O => \N__25999\,
            I => \N__25996\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__25996\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__3760\ : InMux
    port map (
            O => \N__25993\,
            I => \N__25990\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__25990\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25987\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__3757\ : InMux
    port map (
            O => \N__25984\,
            I => \N__25978\
        );

    \I__3756\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25978\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__25978\,
            I => \N__25971\
        );

    \I__3754\ : InMux
    port map (
            O => \N__25977\,
            I => \N__25968\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25961\
        );

    \I__3752\ : InMux
    port map (
            O => \N__25975\,
            I => \N__25961\
        );

    \I__3751\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25961\
        );

    \I__3750\ : Odrv12
    port map (
            O => \N__25971\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__25968\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__25961\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25954\,
            I => \N__25951\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__25951\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__3745\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25945\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__25945\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25942\,
            I => \N__25939\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__25939\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__3741\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25933\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__25933\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__3739\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25927\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__25927\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__3737\ : InMux
    port map (
            O => \N__25924\,
            I => \N__25921\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__25921\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__3735\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25915\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__25915\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__3733\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25909\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__25909\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__25906\,
            I => \N__25903\
        );

    \I__3730\ : InMux
    port map (
            O => \N__25903\,
            I => \N__25900\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__25900\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__3728\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25894\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__25894\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__25891\,
            I => \N__25888\
        );

    \I__3725\ : InMux
    port map (
            O => \N__25888\,
            I => \N__25885\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__25885\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__3723\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25879\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__25879\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__3721\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25873\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__25873\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__3719\ : CascadeMux
    port map (
            O => \N__25870\,
            I => \N__25867\
        );

    \I__3718\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25864\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__25864\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__3716\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25858\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__25858\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__3714\ : CascadeMux
    port map (
            O => \N__25855\,
            I => \N__25852\
        );

    \I__3713\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25849\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__25849\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__3711\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25843\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__25843\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__3709\ : InMux
    port map (
            O => \N__25840\,
            I => \N__25837\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__25837\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__3707\ : InMux
    port map (
            O => \N__25834\,
            I => \N__25831\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__25831\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25825\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__25825\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__3703\ : InMux
    port map (
            O => \N__25822\,
            I => \N__25819\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__25819\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__3701\ : InMux
    port map (
            O => \N__25816\,
            I => \N__25809\
        );

    \I__3700\ : InMux
    port map (
            O => \N__25815\,
            I => \N__25809\
        );

    \I__3699\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25803\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__25809\,
            I => \N__25800\
        );

    \I__3697\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25797\
        );

    \I__3696\ : InMux
    port map (
            O => \N__25807\,
            I => \N__25792\
        );

    \I__3695\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25792\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__25803\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__25800\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__25797\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__25792\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3690\ : InMux
    port map (
            O => \N__25783\,
            I => \N__25779\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__25782\,
            I => \N__25775\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__25779\,
            I => \N__25771\
        );

    \I__3687\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25768\
        );

    \I__3686\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25763\
        );

    \I__3685\ : InMux
    port map (
            O => \N__25774\,
            I => \N__25763\
        );

    \I__3684\ : Span4Mux_h
    port map (
            O => \N__25771\,
            I => \N__25758\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__25768\,
            I => \N__25758\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__25763\,
            I => \N__25755\
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__25758\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__25755\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__3679\ : InMux
    port map (
            O => \N__25750\,
            I => \N__25747\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__25747\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\
        );

    \I__3677\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25741\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__25741\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\
        );

    \I__3675\ : InMux
    port map (
            O => \N__25738\,
            I => \N__25734\
        );

    \I__3674\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25731\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__25734\,
            I => \N__25725\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__25731\,
            I => \N__25725\
        );

    \I__3671\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25722\
        );

    \I__3670\ : Span4Mux_h
    port map (
            O => \N__25725\,
            I => \N__25719\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__25722\,
            I => \N__25714\
        );

    \I__3668\ : Sp12to4
    port map (
            O => \N__25719\,
            I => \N__25714\
        );

    \I__3667\ : Odrv12
    port map (
            O => \N__25714\,
            I => \il_max_comp2_D2\
        );

    \I__3666\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25708\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__25708\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\
        );

    \I__3664\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25701\
        );

    \I__3663\ : InMux
    port map (
            O => \N__25704\,
            I => \N__25698\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__25701\,
            I => \N__25695\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__25698\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__3660\ : Odrv4
    port map (
            O => \N__25695\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__3659\ : CascadeMux
    port map (
            O => \N__25690\,
            I => \N__25687\
        );

    \I__3658\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25684\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__25684\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\
        );

    \I__3656\ : CascadeMux
    port map (
            O => \N__25681\,
            I => \N__25677\
        );

    \I__3655\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25674\
        );

    \I__3654\ : InMux
    port map (
            O => \N__25677\,
            I => \N__25671\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__25674\,
            I => \N__25668\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__25671\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__3651\ : Odrv4
    port map (
            O => \N__25668\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__3650\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25645\
        );

    \I__3649\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25645\
        );

    \I__3648\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25645\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__25660\,
            I => \N__25634\
        );

    \I__3646\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25626\
        );

    \I__3645\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25626\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25657\,
            I => \N__25613\
        );

    \I__3643\ : InMux
    port map (
            O => \N__25656\,
            I => \N__25613\
        );

    \I__3642\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25613\
        );

    \I__3641\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25613\
        );

    \I__3640\ : InMux
    port map (
            O => \N__25653\,
            I => \N__25613\
        );

    \I__3639\ : InMux
    port map (
            O => \N__25652\,
            I => \N__25613\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__25645\,
            I => \N__25610\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25644\,
            I => \N__25593\
        );

    \I__3636\ : InMux
    port map (
            O => \N__25643\,
            I => \N__25593\
        );

    \I__3635\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25593\
        );

    \I__3634\ : InMux
    port map (
            O => \N__25641\,
            I => \N__25593\
        );

    \I__3633\ : InMux
    port map (
            O => \N__25640\,
            I => \N__25593\
        );

    \I__3632\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25593\
        );

    \I__3631\ : InMux
    port map (
            O => \N__25638\,
            I => \N__25593\
        );

    \I__3630\ : InMux
    port map (
            O => \N__25637\,
            I => \N__25593\
        );

    \I__3629\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25588\
        );

    \I__3628\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25588\
        );

    \I__3627\ : InMux
    port map (
            O => \N__25632\,
            I => \N__25582\
        );

    \I__3626\ : InMux
    port map (
            O => \N__25631\,
            I => \N__25582\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__25626\,
            I => \N__25577\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__25613\,
            I => \N__25577\
        );

    \I__3623\ : Span4Mux_v
    port map (
            O => \N__25610\,
            I => \N__25574\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__25593\,
            I => \N__25569\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__25588\,
            I => \N__25569\
        );

    \I__3620\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25566\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__25582\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__25577\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__25574\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3616\ : Odrv12
    port map (
            O => \N__25569\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__25566\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__25555\,
            I => \N__25544\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__25554\,
            I => \N__25541\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__25553\,
            I => \N__25538\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__25552\,
            I => \N__25535\
        );

    \I__3610\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25524\
        );

    \I__3609\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25524\
        );

    \I__3608\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25517\
        );

    \I__3607\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25517\
        );

    \I__3606\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25517\
        );

    \I__3605\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25500\
        );

    \I__3604\ : InMux
    port map (
            O => \N__25541\,
            I => \N__25500\
        );

    \I__3603\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25500\
        );

    \I__3602\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25500\
        );

    \I__3601\ : InMux
    port map (
            O => \N__25534\,
            I => \N__25487\
        );

    \I__3600\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25487\
        );

    \I__3599\ : InMux
    port map (
            O => \N__25532\,
            I => \N__25487\
        );

    \I__3598\ : InMux
    port map (
            O => \N__25531\,
            I => \N__25487\
        );

    \I__3597\ : InMux
    port map (
            O => \N__25530\,
            I => \N__25487\
        );

    \I__3596\ : InMux
    port map (
            O => \N__25529\,
            I => \N__25487\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__25524\,
            I => \N__25482\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__25517\,
            I => \N__25482\
        );

    \I__3593\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25477\
        );

    \I__3592\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25477\
        );

    \I__3591\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25471\
        );

    \I__3590\ : InMux
    port map (
            O => \N__25513\,
            I => \N__25471\
        );

    \I__3589\ : InMux
    port map (
            O => \N__25512\,
            I => \N__25462\
        );

    \I__3588\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25462\
        );

    \I__3587\ : InMux
    port map (
            O => \N__25510\,
            I => \N__25462\
        );

    \I__3586\ : InMux
    port map (
            O => \N__25509\,
            I => \N__25462\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__25500\,
            I => \N__25455\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__25487\,
            I => \N__25455\
        );

    \I__3583\ : Span4Mux_h
    port map (
            O => \N__25482\,
            I => \N__25455\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__25477\,
            I => \N__25452\
        );

    \I__3581\ : InMux
    port map (
            O => \N__25476\,
            I => \N__25449\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__25471\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__25462\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__25455\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3577\ : Odrv12
    port map (
            O => \N__25452\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__25449\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__25438\,
            I => \N__25424\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__25437\,
            I => \N__25421\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__25436\,
            I => \N__25414\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__25435\,
            I => \N__25411\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__25434\,
            I => \N__25408\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__25433\,
            I => \N__25405\
        );

    \I__3569\ : CascadeMux
    port map (
            O => \N__25432\,
            I => \N__25402\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__25431\,
            I => \N__25399\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__25430\,
            I => \N__25396\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__25429\,
            I => \N__25393\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__25428\,
            I => \N__25390\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__25427\,
            I => \N__25382\
        );

    \I__3563\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25375\
        );

    \I__3562\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25375\
        );

    \I__3561\ : InMux
    port map (
            O => \N__25420\,
            I => \N__25375\
        );

    \I__3560\ : InMux
    port map (
            O => \N__25419\,
            I => \N__25360\
        );

    \I__3559\ : InMux
    port map (
            O => \N__25418\,
            I => \N__25360\
        );

    \I__3558\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25360\
        );

    \I__3557\ : InMux
    port map (
            O => \N__25414\,
            I => \N__25360\
        );

    \I__3556\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25360\
        );

    \I__3555\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25360\
        );

    \I__3554\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25355\
        );

    \I__3553\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25355\
        );

    \I__3552\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25338\
        );

    \I__3551\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25338\
        );

    \I__3550\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25338\
        );

    \I__3549\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25338\
        );

    \I__3548\ : InMux
    port map (
            O => \N__25389\,
            I => \N__25338\
        );

    \I__3547\ : InMux
    port map (
            O => \N__25388\,
            I => \N__25338\
        );

    \I__3546\ : InMux
    port map (
            O => \N__25387\,
            I => \N__25338\
        );

    \I__3545\ : InMux
    port map (
            O => \N__25386\,
            I => \N__25338\
        );

    \I__3544\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25333\
        );

    \I__3543\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25333\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__25375\,
            I => \N__25330\
        );

    \I__3541\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25325\
        );

    \I__3540\ : InMux
    port map (
            O => \N__25373\,
            I => \N__25325\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__25360\,
            I => \N__25321\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__25355\,
            I => \N__25314\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__25338\,
            I => \N__25314\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__25333\,
            I => \N__25314\
        );

    \I__3535\ : Span4Mux_v
    port map (
            O => \N__25330\,
            I => \N__25309\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__25325\,
            I => \N__25309\
        );

    \I__3533\ : InMux
    port map (
            O => \N__25324\,
            I => \N__25306\
        );

    \I__3532\ : Span4Mux_v
    port map (
            O => \N__25321\,
            I => \N__25301\
        );

    \I__3531\ : Span4Mux_v
    port map (
            O => \N__25314\,
            I => \N__25301\
        );

    \I__3530\ : Span4Mux_h
    port map (
            O => \N__25309\,
            I => \N__25298\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__25306\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3528\ : Odrv4
    port map (
            O => \N__25301\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3527\ : Odrv4
    port map (
            O => \N__25298\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__3526\ : InMux
    port map (
            O => \N__25291\,
            I => \N__25288\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__25288\,
            I => \N__25285\
        );

    \I__3524\ : Odrv4
    port map (
            O => \N__25285\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__25282\,
            I => \N__25279\
        );

    \I__3522\ : InMux
    port map (
            O => \N__25279\,
            I => \N__25276\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__25276\,
            I => \N__25272\
        );

    \I__3520\ : InMux
    port map (
            O => \N__25275\,
            I => \N__25269\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__25272\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__25269\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__25264\,
            I => \N__25261\
        );

    \I__3516\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25258\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__25258\,
            I => \N__25255\
        );

    \I__3514\ : Span4Mux_h
    port map (
            O => \N__25255\,
            I => \N__25252\
        );

    \I__3513\ : Odrv4
    port map (
            O => \N__25252\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__25249\,
            I => \N__25246\
        );

    \I__3511\ : InMux
    port map (
            O => \N__25246\,
            I => \N__25243\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__25243\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__25240\,
            I => \N__25237\
        );

    \I__3508\ : InMux
    port map (
            O => \N__25237\,
            I => \N__25234\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__25234\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__25231\,
            I => \N__25228\
        );

    \I__3505\ : InMux
    port map (
            O => \N__25228\,
            I => \N__25225\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__25225\,
            I => \N__25222\
        );

    \I__3503\ : Odrv12
    port map (
            O => \N__25222\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__25219\,
            I => \N__25216\
        );

    \I__3501\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25213\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__25213\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__25210\,
            I => \N__25207\
        );

    \I__3498\ : InMux
    port map (
            O => \N__25207\,
            I => \N__25204\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__25204\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__25201\,
            I => \N__25198\
        );

    \I__3495\ : InMux
    port map (
            O => \N__25198\,
            I => \N__25195\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__25195\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__3493\ : CEMux
    port map (
            O => \N__25192\,
            I => \N__25186\
        );

    \I__3492\ : CEMux
    port map (
            O => \N__25191\,
            I => \N__25183\
        );

    \I__3491\ : CEMux
    port map (
            O => \N__25190\,
            I => \N__25180\
        );

    \I__3490\ : CEMux
    port map (
            O => \N__25189\,
            I => \N__25177\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__25186\,
            I => \N__25173\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__25183\,
            I => \N__25170\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__25180\,
            I => \N__25167\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25164\
        );

    \I__3485\ : CEMux
    port map (
            O => \N__25176\,
            I => \N__25161\
        );

    \I__3484\ : Span4Mux_v
    port map (
            O => \N__25173\,
            I => \N__25158\
        );

    \I__3483\ : Span4Mux_h
    port map (
            O => \N__25170\,
            I => \N__25155\
        );

    \I__3482\ : Span4Mux_v
    port map (
            O => \N__25167\,
            I => \N__25152\
        );

    \I__3481\ : Span4Mux_h
    port map (
            O => \N__25164\,
            I => \N__25147\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__25161\,
            I => \N__25147\
        );

    \I__3479\ : Odrv4
    port map (
            O => \N__25158\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__25155\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__25152\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__3476\ : Odrv4
    port map (
            O => \N__25147\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__25138\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_\
        );

    \I__3474\ : InMux
    port map (
            O => \N__25135\,
            I => \N__25129\
        );

    \I__3473\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25126\
        );

    \I__3472\ : InMux
    port map (
            O => \N__25133\,
            I => \N__25123\
        );

    \I__3471\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25120\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__25129\,
            I => \N__25117\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__25126\,
            I => \N__25114\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__25123\,
            I => \N__25111\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__25120\,
            I => \N__25104\
        );

    \I__3466\ : Span4Mux_h
    port map (
            O => \N__25117\,
            I => \N__25104\
        );

    \I__3465\ : Span4Mux_h
    port map (
            O => \N__25114\,
            I => \N__25099\
        );

    \I__3464\ : Span4Mux_h
    port map (
            O => \N__25111\,
            I => \N__25099\
        );

    \I__3463\ : InMux
    port map (
            O => \N__25110\,
            I => \N__25096\
        );

    \I__3462\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25093\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__25104\,
            I => phase_controller_inst1_state_4
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__25099\,
            I => phase_controller_inst1_state_4
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__25096\,
            I => phase_controller_inst1_state_4
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__25093\,
            I => phase_controller_inst1_state_4
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__25084\,
            I => \N__25081\
        );

    \I__3456\ : InMux
    port map (
            O => \N__25081\,
            I => \N__25078\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__25078\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__25075\,
            I => \N__25072\
        );

    \I__3453\ : InMux
    port map (
            O => \N__25072\,
            I => \N__25069\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__25069\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__25066\,
            I => \N__25063\
        );

    \I__3450\ : InMux
    port map (
            O => \N__25063\,
            I => \N__25060\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__25060\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__25057\,
            I => \N__25054\
        );

    \I__3447\ : InMux
    port map (
            O => \N__25054\,
            I => \N__25051\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__25051\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__3445\ : CascadeMux
    port map (
            O => \N__25048\,
            I => \N__25045\
        );

    \I__3444\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25042\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__25042\,
            I => \N__25039\
        );

    \I__3442\ : Span4Mux_v
    port map (
            O => \N__25039\,
            I => \N__25036\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__25036\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__3440\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25030\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__25030\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__25027\,
            I => \N__25024\
        );

    \I__3437\ : InMux
    port map (
            O => \N__25024\,
            I => \N__25021\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__25021\,
            I => \N__25018\
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__25018\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__25015\,
            I => \N__25012\
        );

    \I__3433\ : InMux
    port map (
            O => \N__25012\,
            I => \N__25009\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__25009\,
            I => \N__25006\
        );

    \I__3431\ : Span4Mux_v
    port map (
            O => \N__25006\,
            I => \N__25003\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__25003\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__3429\ : CascadeMux
    port map (
            O => \N__25000\,
            I => \N__24997\
        );

    \I__3428\ : InMux
    port map (
            O => \N__24997\,
            I => \N__24994\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__24994\,
            I => \N__24991\
        );

    \I__3426\ : Span4Mux_h
    port map (
            O => \N__24991\,
            I => \N__24988\
        );

    \I__3425\ : Odrv4
    port map (
            O => \N__24988\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__3424\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24981\
        );

    \I__3423\ : InMux
    port map (
            O => \N__24984\,
            I => \N__24978\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__24981\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__24978\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__3420\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24970\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__24970\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__3418\ : InMux
    port map (
            O => \N__24967\,
            I => \N__24963\
        );

    \I__3417\ : InMux
    port map (
            O => \N__24966\,
            I => \N__24960\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__24963\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__24960\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__3414\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24952\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__24952\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__3412\ : InMux
    port map (
            O => \N__24949\,
            I => \N__24945\
        );

    \I__3411\ : InMux
    port map (
            O => \N__24948\,
            I => \N__24942\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__24945\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__24942\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24934\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__24934\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__3406\ : InMux
    port map (
            O => \N__24931\,
            I => \N__24928\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__24928\,
            I => \N__24924\
        );

    \I__3404\ : InMux
    port map (
            O => \N__24927\,
            I => \N__24921\
        );

    \I__3403\ : Span4Mux_h
    port map (
            O => \N__24924\,
            I => \N__24918\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__24921\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__24918\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__3400\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24910\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__24910\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\
        );

    \I__3398\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24903\
        );

    \I__3397\ : InMux
    port map (
            O => \N__24906\,
            I => \N__24900\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__24903\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__24900\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__3394\ : InMux
    port map (
            O => \N__24895\,
            I => \N__24892\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__24892\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\
        );

    \I__3392\ : InMux
    port map (
            O => \N__24889\,
            I => \N__24885\
        );

    \I__3391\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24882\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__24885\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__24882\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__3388\ : InMux
    port map (
            O => \N__24877\,
            I => \N__24874\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__24874\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\
        );

    \I__3386\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24867\
        );

    \I__3385\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24864\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__24867\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__24864\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__3382\ : InMux
    port map (
            O => \N__24859\,
            I => \N__24856\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__24856\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\
        );

    \I__3380\ : InMux
    port map (
            O => \N__24853\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__3379\ : InMux
    port map (
            O => \N__24850\,
            I => \N__24847\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__24847\,
            I => \N__24843\
        );

    \I__3377\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24840\
        );

    \I__3376\ : Odrv4
    port map (
            O => \N__24843\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__24840\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__3374\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24832\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__24832\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__24829\,
            I => \N__24826\
        );

    \I__3371\ : InMux
    port map (
            O => \N__24826\,
            I => \N__24823\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__24823\,
            I => \N__24820\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__24820\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__24817\,
            I => \N__24814\
        );

    \I__3367\ : InMux
    port map (
            O => \N__24814\,
            I => \N__24811\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__24811\,
            I => \N__24807\
        );

    \I__3365\ : InMux
    port map (
            O => \N__24810\,
            I => \N__24804\
        );

    \I__3364\ : Odrv4
    port map (
            O => \N__24807\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__24804\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__3362\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24796\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__24796\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__24793\,
            I => \N__24790\
        );

    \I__3359\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24787\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__24787\,
            I => \N__24783\
        );

    \I__3357\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24780\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__24783\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__24780\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__3354\ : InMux
    port map (
            O => \N__24775\,
            I => \N__24772\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__24772\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__24769\,
            I => \N__24766\
        );

    \I__3351\ : InMux
    port map (
            O => \N__24766\,
            I => \N__24763\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__24763\,
            I => \N__24759\
        );

    \I__3349\ : InMux
    port map (
            O => \N__24762\,
            I => \N__24756\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__24759\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__24756\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__3346\ : InMux
    port map (
            O => \N__24751\,
            I => \N__24748\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__24748\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__3344\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24741\
        );

    \I__3343\ : InMux
    port map (
            O => \N__24744\,
            I => \N__24738\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__24741\,
            I => \N__24735\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__24738\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__24735\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__3339\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24727\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__24727\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__3337\ : InMux
    port map (
            O => \N__24724\,
            I => \N__24720\
        );

    \I__3336\ : InMux
    port map (
            O => \N__24723\,
            I => \N__24717\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__24720\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__24717\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__3333\ : InMux
    port map (
            O => \N__24712\,
            I => \N__24709\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__24709\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__3331\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24702\
        );

    \I__3330\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24699\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__24702\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__24699\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__3327\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24691\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__24691\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__3325\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24684\
        );

    \I__3324\ : InMux
    port map (
            O => \N__24687\,
            I => \N__24681\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__24684\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__24681\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__3321\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24673\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__24673\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__3319\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24666\
        );

    \I__3318\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24663\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__24666\,
            I => \N__24658\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__24663\,
            I => \N__24658\
        );

    \I__3315\ : Span4Mux_v
    port map (
            O => \N__24658\,
            I => \N__24655\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__24655\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__3313\ : InMux
    port map (
            O => \N__24652\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__3312\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24646\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24642\
        );

    \I__3310\ : InMux
    port map (
            O => \N__24645\,
            I => \N__24639\
        );

    \I__3309\ : Span4Mux_v
    port map (
            O => \N__24642\,
            I => \N__24634\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__24639\,
            I => \N__24634\
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__24634\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__3306\ : InMux
    port map (
            O => \N__24631\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__3305\ : InMux
    port map (
            O => \N__24628\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__24625\,
            I => \N__24621\
        );

    \I__3303\ : CascadeMux
    port map (
            O => \N__24624\,
            I => \N__24618\
        );

    \I__3302\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24609\
        );

    \I__3301\ : InMux
    port map (
            O => \N__24618\,
            I => \N__24609\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__24617\,
            I => \N__24605\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__24616\,
            I => \N__24602\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__24615\,
            I => \N__24597\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__24614\,
            I => \N__24594\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__24609\,
            I => \N__24590\
        );

    \I__3295\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24581\
        );

    \I__3294\ : InMux
    port map (
            O => \N__24605\,
            I => \N__24581\
        );

    \I__3293\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24581\
        );

    \I__3292\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24581\
        );

    \I__3291\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24578\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24597\,
            I => \N__24575\
        );

    \I__3289\ : InMux
    port map (
            O => \N__24594\,
            I => \N__24570\
        );

    \I__3288\ : InMux
    port map (
            O => \N__24593\,
            I => \N__24570\
        );

    \I__3287\ : Span4Mux_v
    port map (
            O => \N__24590\,
            I => \N__24563\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__24581\,
            I => \N__24563\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__24578\,
            I => \N__24563\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__24575\,
            I => \N__24558\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__24570\,
            I => \N__24558\
        );

    \I__3282\ : Span4Mux_h
    port map (
            O => \N__24563\,
            I => \N__24555\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__24558\,
            I => \N__24552\
        );

    \I__3280\ : Span4Mux_v
    port map (
            O => \N__24555\,
            I => \N__24549\
        );

    \I__3279\ : Span4Mux_v
    port map (
            O => \N__24552\,
            I => \N__24546\
        );

    \I__3278\ : Span4Mux_h
    port map (
            O => \N__24549\,
            I => \N__24543\
        );

    \I__3277\ : Span4Mux_h
    port map (
            O => \N__24546\,
            I => \N__24540\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__24543\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__24540\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__24535\,
            I => \N__24531\
        );

    \I__3273\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24528\
        );

    \I__3272\ : InMux
    port map (
            O => \N__24531\,
            I => \N__24525\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__24528\,
            I => \N__24519\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__24525\,
            I => \N__24519\
        );

    \I__3269\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24516\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__24519\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__24516\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__3266\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24508\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__24508\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__3264\ : InMux
    port map (
            O => \N__24505\,
            I => \N__24502\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__24502\,
            I => \N__24498\
        );

    \I__3262\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24495\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__24498\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__24495\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__3259\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24487\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__24487\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__24484\,
            I => \N__24481\
        );

    \I__3256\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24478\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__24478\,
            I => \N__24474\
        );

    \I__3254\ : InMux
    port map (
            O => \N__24477\,
            I => \N__24471\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__24474\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__24471\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__3251\ : InMux
    port map (
            O => \N__24466\,
            I => \N__24463\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__24463\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__3249\ : InMux
    port map (
            O => \N__24460\,
            I => \N__24456\
        );

    \I__3248\ : InMux
    port map (
            O => \N__24459\,
            I => \N__24453\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24450\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__24453\,
            I => \N__24447\
        );

    \I__3245\ : Odrv4
    port map (
            O => \N__24450\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__24447\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__3243\ : InMux
    port map (
            O => \N__24442\,
            I => \N__24439\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__24439\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__3241\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24430\
        );

    \I__3240\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24430\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__24430\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__3238\ : InMux
    port map (
            O => \N__24427\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__3237\ : InMux
    port map (
            O => \N__24424\,
            I => \N__24420\
        );

    \I__3236\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24417\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__24420\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__24417\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__3233\ : InMux
    port map (
            O => \N__24412\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__3232\ : CascadeMux
    port map (
            O => \N__24409\,
            I => \N__24405\
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__24408\,
            I => \N__24402\
        );

    \I__3230\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24397\
        );

    \I__3229\ : InMux
    port map (
            O => \N__24402\,
            I => \N__24397\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__24397\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__3227\ : InMux
    port map (
            O => \N__24394\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__3226\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24385\
        );

    \I__3225\ : InMux
    port map (
            O => \N__24390\,
            I => \N__24385\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__24385\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__3223\ : InMux
    port map (
            O => \N__24382\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__3222\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24376\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__24376\,
            I => \N__24372\
        );

    \I__3220\ : InMux
    port map (
            O => \N__24375\,
            I => \N__24369\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__24372\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__24369\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__3217\ : InMux
    port map (
            O => \N__24364\,
            I => \bfn_9_11_0_\
        );

    \I__3216\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24357\
        );

    \I__3215\ : InMux
    port map (
            O => \N__24360\,
            I => \N__24354\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__24357\,
            I => \N__24351\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__24354\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__24351\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__3211\ : InMux
    port map (
            O => \N__24346\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__3210\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24339\
        );

    \I__3209\ : InMux
    port map (
            O => \N__24342\,
            I => \N__24336\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__24339\,
            I => \N__24333\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__24336\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__3206\ : Odrv4
    port map (
            O => \N__24333\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__3205\ : InMux
    port map (
            O => \N__24328\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__24325\,
            I => \N__24321\
        );

    \I__3203\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24318\
        );

    \I__3202\ : InMux
    port map (
            O => \N__24321\,
            I => \N__24315\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__24318\,
            I => \N__24312\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__24315\,
            I => \N__24309\
        );

    \I__3199\ : Odrv4
    port map (
            O => \N__24312\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__24309\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__3197\ : InMux
    port map (
            O => \N__24304\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__3196\ : InMux
    port map (
            O => \N__24301\,
            I => \N__24298\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__24298\,
            I => \N__24294\
        );

    \I__3194\ : InMux
    port map (
            O => \N__24297\,
            I => \N__24291\
        );

    \I__3193\ : Span4Mux_v
    port map (
            O => \N__24294\,
            I => \N__24288\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__24291\,
            I => \N__24285\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__24288\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__24285\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__3189\ : InMux
    port map (
            O => \N__24280\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__3188\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24271\
        );

    \I__3187\ : InMux
    port map (
            O => \N__24276\,
            I => \N__24271\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__24271\,
            I => \N__24268\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__24268\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__3184\ : InMux
    port map (
            O => \N__24265\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__3183\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24256\
        );

    \I__3182\ : InMux
    port map (
            O => \N__24261\,
            I => \N__24256\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__24256\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__3180\ : InMux
    port map (
            O => \N__24253\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__24250\,
            I => \N__24247\
        );

    \I__3178\ : InMux
    port map (
            O => \N__24247\,
            I => \N__24244\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__24244\,
            I => \N__24241\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__24241\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__3175\ : CascadeMux
    port map (
            O => \N__24238\,
            I => \N__24235\
        );

    \I__3174\ : InMux
    port map (
            O => \N__24235\,
            I => \N__24229\
        );

    \I__3173\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24229\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__24229\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__3171\ : InMux
    port map (
            O => \N__24226\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__3170\ : InMux
    port map (
            O => \N__24223\,
            I => \N__24219\
        );

    \I__3169\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24216\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__24219\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__24216\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__3166\ : InMux
    port map (
            O => \N__24211\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__3165\ : InMux
    port map (
            O => \N__24208\,
            I => \N__24204\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__24207\,
            I => \N__24201\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__24204\,
            I => \N__24198\
        );

    \I__3162\ : InMux
    port map (
            O => \N__24201\,
            I => \N__24195\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__24198\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__24195\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__3159\ : InMux
    port map (
            O => \N__24190\,
            I => \bfn_9_10_0_\
        );

    \I__3158\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24183\
        );

    \I__3157\ : InMux
    port map (
            O => \N__24186\,
            I => \N__24180\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__24183\,
            I => \N__24177\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__24180\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__24177\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__3153\ : InMux
    port map (
            O => \N__24172\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__24169\,
            I => \N__24166\
        );

    \I__3151\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24162\
        );

    \I__3150\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24159\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__24162\,
            I => \N__24156\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__24159\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__3147\ : Odrv4
    port map (
            O => \N__24156\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__3146\ : InMux
    port map (
            O => \N__24151\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__3145\ : InMux
    port map (
            O => \N__24148\,
            I => \N__24142\
        );

    \I__3144\ : InMux
    port map (
            O => \N__24147\,
            I => \N__24142\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__24142\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__3142\ : InMux
    port map (
            O => \N__24139\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__3141\ : InMux
    port map (
            O => \N__24136\,
            I => \N__24132\
        );

    \I__3140\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24127\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__24132\,
            I => \N__24124\
        );

    \I__3138\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24121\
        );

    \I__3137\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24118\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__24127\,
            I => \N__24115\
        );

    \I__3135\ : Span4Mux_v
    port map (
            O => \N__24124\,
            I => \N__24110\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__24121\,
            I => \N__24110\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__24118\,
            I => \N__24107\
        );

    \I__3132\ : Span4Mux_v
    port map (
            O => \N__24115\,
            I => \N__24104\
        );

    \I__3131\ : Span4Mux_h
    port map (
            O => \N__24110\,
            I => \N__24101\
        );

    \I__3130\ : Span12Mux_s7_v
    port map (
            O => \N__24107\,
            I => \N__24098\
        );

    \I__3129\ : Span4Mux_h
    port map (
            O => \N__24104\,
            I => \N__24095\
        );

    \I__3128\ : Span4Mux_h
    port map (
            O => \N__24101\,
            I => \N__24092\
        );

    \I__3127\ : Odrv12
    port map (
            O => \N__24098\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__24095\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__24092\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__3124\ : InMux
    port map (
            O => \N__24085\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__3123\ : InMux
    port map (
            O => \N__24082\,
            I => \N__24079\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__24079\,
            I => \N__24074\
        );

    \I__3121\ : InMux
    port map (
            O => \N__24078\,
            I => \N__24071\
        );

    \I__3120\ : InMux
    port map (
            O => \N__24077\,
            I => \N__24068\
        );

    \I__3119\ : Span4Mux_v
    port map (
            O => \N__24074\,
            I => \N__24061\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__24071\,
            I => \N__24061\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__24068\,
            I => \N__24061\
        );

    \I__3116\ : Span4Mux_h
    port map (
            O => \N__24061\,
            I => \N__24058\
        );

    \I__3115\ : Span4Mux_h
    port map (
            O => \N__24058\,
            I => \N__24055\
        );

    \I__3114\ : Odrv4
    port map (
            O => \N__24055\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__3113\ : InMux
    port map (
            O => \N__24052\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__3112\ : InMux
    port map (
            O => \N__24049\,
            I => \N__24044\
        );

    \I__3111\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24041\
        );

    \I__3110\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24038\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__24044\,
            I => \N__24031\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__24041\,
            I => \N__24031\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__24038\,
            I => \N__24031\
        );

    \I__3106\ : Span4Mux_h
    port map (
            O => \N__24031\,
            I => \N__24028\
        );

    \I__3105\ : Span4Mux_h
    port map (
            O => \N__24028\,
            I => \N__24025\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__24025\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__3103\ : InMux
    port map (
            O => \N__24022\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__3102\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24014\
        );

    \I__3101\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24011\
        );

    \I__3100\ : InMux
    port map (
            O => \N__24017\,
            I => \N__24008\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__24014\,
            I => \N__24001\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__24001\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__24008\,
            I => \N__24001\
        );

    \I__3096\ : Span4Mux_h
    port map (
            O => \N__24001\,
            I => \N__23998\
        );

    \I__3095\ : Span4Mux_h
    port map (
            O => \N__23998\,
            I => \N__23995\
        );

    \I__3094\ : Odrv4
    port map (
            O => \N__23995\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23992\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__3092\ : InMux
    port map (
            O => \N__23989\,
            I => \N__23986\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23986\,
            I => \N__23981\
        );

    \I__3090\ : InMux
    port map (
            O => \N__23985\,
            I => \N__23978\
        );

    \I__3089\ : InMux
    port map (
            O => \N__23984\,
            I => \N__23975\
        );

    \I__3088\ : Span4Mux_v
    port map (
            O => \N__23981\,
            I => \N__23968\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__23978\,
            I => \N__23968\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__23975\,
            I => \N__23968\
        );

    \I__3085\ : Span4Mux_h
    port map (
            O => \N__23968\,
            I => \N__23965\
        );

    \I__3084\ : Span4Mux_h
    port map (
            O => \N__23965\,
            I => \N__23962\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__23962\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__3082\ : InMux
    port map (
            O => \N__23959\,
            I => \bfn_9_9_0_\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23952\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23949\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__23952\,
            I => \N__23943\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__23949\,
            I => \N__23943\
        );

    \I__3077\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23940\
        );

    \I__3076\ : Sp12to4
    port map (
            O => \N__23943\,
            I => \N__23935\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__23940\,
            I => \N__23935\
        );

    \I__3074\ : Span12Mux_s9_h
    port map (
            O => \N__23935\,
            I => \N__23932\
        );

    \I__3073\ : Odrv12
    port map (
            O => \N__23932\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__3072\ : InMux
    port map (
            O => \N__23929\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__23926\,
            I => \N__23923\
        );

    \I__3070\ : InMux
    port map (
            O => \N__23923\,
            I => \N__23920\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__23920\,
            I => \N__23916\
        );

    \I__3068\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23913\
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__23916\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__23913\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__3065\ : InMux
    port map (
            O => \N__23908\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__3064\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23899\
        );

    \I__3063\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23899\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__23899\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__3061\ : InMux
    port map (
            O => \N__23896\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__3060\ : CascadeMux
    port map (
            O => \N__23893\,
            I => \N__23890\
        );

    \I__3059\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23887\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__23887\,
            I => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__3057\ : InMux
    port map (
            O => \N__23884\,
            I => \N__23881\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__23881\,
            I => \N__23877\
        );

    \I__3055\ : InMux
    port map (
            O => \N__23880\,
            I => \N__23874\
        );

    \I__3054\ : Span4Mux_v
    port map (
            O => \N__23877\,
            I => \N__23868\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__23874\,
            I => \N__23868\
        );

    \I__3052\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23865\
        );

    \I__3051\ : Span4Mux_h
    port map (
            O => \N__23868\,
            I => \N__23859\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__23865\,
            I => \N__23859\
        );

    \I__3049\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23856\
        );

    \I__3048\ : Sp12to4
    port map (
            O => \N__23859\,
            I => \N__23853\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__23856\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__3046\ : Odrv12
    port map (
            O => \N__23853\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__3045\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23845\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__23845\,
            I => \N__23842\
        );

    \I__3043\ : Glb2LocalMux
    port map (
            O => \N__23842\,
            I => \N__23839\
        );

    \I__3042\ : GlobalMux
    port map (
            O => \N__23839\,
            I => clk_12mhz
        );

    \I__3041\ : IoInMux
    port map (
            O => \N__23836\,
            I => \N__23833\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__23833\,
            I => \N__23830\
        );

    \I__3039\ : Span4Mux_s0_v
    port map (
            O => \N__23830\,
            I => \N__23827\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__23827\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__3037\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23821\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__23821\,
            I => \N__23818\
        );

    \I__3035\ : Odrv12
    port map (
            O => \N__23818\,
            I => il_min_comp1_c
        );

    \I__3034\ : InMux
    port map (
            O => \N__23815\,
            I => \N__23812\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__23812\,
            I => \N__23809\
        );

    \I__3032\ : Span4Mux_h
    port map (
            O => \N__23809\,
            I => \N__23806\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__23806\,
            I => \il_min_comp1_D1\
        );

    \I__3030\ : InMux
    port map (
            O => \N__23803\,
            I => \N__23800\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__23800\,
            I => \N__23797\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__23797\,
            I => \N__23794\
        );

    \I__3027\ : Span4Mux_h
    port map (
            O => \N__23794\,
            I => \N__23791\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__23791\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__3025\ : InMux
    port map (
            O => \N__23788\,
            I => \N__23785\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__23785\,
            I => \N__23782\
        );

    \I__3023\ : Span12Mux_s9_h
    port map (
            O => \N__23782\,
            I => \N__23779\
        );

    \I__3022\ : Odrv12
    port map (
            O => \N__23779\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__3021\ : InMux
    port map (
            O => \N__23776\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__3020\ : InMux
    port map (
            O => \N__23773\,
            I => \N__23770\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__23770\,
            I => \N__23767\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__23767\,
            I => \N__23764\
        );

    \I__3017\ : Span4Mux_h
    port map (
            O => \N__23764\,
            I => \N__23761\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__23761\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__3015\ : InMux
    port map (
            O => \N__23758\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__3014\ : InMux
    port map (
            O => \N__23755\,
            I => \N__23752\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__23752\,
            I => \N__23748\
        );

    \I__3012\ : InMux
    port map (
            O => \N__23751\,
            I => \N__23745\
        );

    \I__3011\ : Span4Mux_s2_h
    port map (
            O => \N__23748\,
            I => \N__23739\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__23745\,
            I => \N__23739\
        );

    \I__3009\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23736\
        );

    \I__3008\ : Sp12to4
    port map (
            O => \N__23739\,
            I => \N__23731\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__23736\,
            I => \N__23731\
        );

    \I__3006\ : Span12Mux_s7_v
    port map (
            O => \N__23731\,
            I => \N__23728\
        );

    \I__3005\ : Odrv12
    port map (
            O => \N__23728\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__3004\ : InMux
    port map (
            O => \N__23725\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__3003\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23718\
        );

    \I__3002\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23715\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__23718\,
            I => \N__23712\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__23715\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__2999\ : Odrv4
    port map (
            O => \N__23712\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__2998\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23704\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__23704\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\
        );

    \I__2996\ : InMux
    port map (
            O => \N__23701\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__2995\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23694\
        );

    \I__2994\ : InMux
    port map (
            O => \N__23697\,
            I => \N__23691\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__23694\,
            I => \N__23688\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__23691\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__23688\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__23683\,
            I => \N__23680\
        );

    \I__2989\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23677\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__23677\,
            I => \N__23674\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__23674\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\
        );

    \I__2986\ : InMux
    port map (
            O => \N__23671\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__2985\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23665\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__23665\,
            I => \N__23661\
        );

    \I__2983\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23658\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__23661\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__23658\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__23653\,
            I => \N__23650\
        );

    \I__2979\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23647\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__23647\,
            I => \N__23644\
        );

    \I__2977\ : Span4Mux_h
    port map (
            O => \N__23644\,
            I => \N__23641\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__23641\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\
        );

    \I__2975\ : InMux
    port map (
            O => \N__23638\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__2974\ : InMux
    port map (
            O => \N__23635\,
            I => \N__23631\
        );

    \I__2973\ : InMux
    port map (
            O => \N__23634\,
            I => \N__23628\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__23631\,
            I => \N__23625\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__23628\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__23625\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__2969\ : InMux
    port map (
            O => \N__23620\,
            I => \N__23617\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__23617\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\
        );

    \I__2967\ : InMux
    port map (
            O => \N__23614\,
            I => \bfn_8_22_0_\
        );

    \I__2966\ : InMux
    port map (
            O => \N__23611\,
            I => \N__23607\
        );

    \I__2965\ : InMux
    port map (
            O => \N__23610\,
            I => \N__23604\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__23607\,
            I => \N__23601\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__23604\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__2962\ : Odrv4
    port map (
            O => \N__23601\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__2961\ : InMux
    port map (
            O => \N__23596\,
            I => \N__23593\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__23593\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\
        );

    \I__2959\ : InMux
    port map (
            O => \N__23590\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__2958\ : InMux
    port map (
            O => \N__23587\,
            I => \N__23583\
        );

    \I__2957\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23580\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__23583\,
            I => \N__23577\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__23580\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__23577\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__2953\ : InMux
    port map (
            O => \N__23572\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__2952\ : InMux
    port map (
            O => \N__23569\,
            I => \N__23566\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__23566\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\
        );

    \I__2950\ : InMux
    port map (
            O => \N__23563\,
            I => \N__23560\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__23560\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\
        );

    \I__2948\ : InMux
    port map (
            O => \N__23557\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__2947\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23550\
        );

    \I__2946\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23547\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__23550\,
            I => \N__23542\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__23547\,
            I => \N__23542\
        );

    \I__2943\ : Span4Mux_v
    port map (
            O => \N__23542\,
            I => \N__23539\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__23539\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__2941\ : InMux
    port map (
            O => \N__23536\,
            I => \N__23533\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__23533\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\
        );

    \I__2939\ : InMux
    port map (
            O => \N__23530\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__2938\ : InMux
    port map (
            O => \N__23527\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__2937\ : InMux
    port map (
            O => \N__23524\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__2936\ : InMux
    port map (
            O => \N__23521\,
            I => \bfn_8_21_0_\
        );

    \I__2935\ : InMux
    port map (
            O => \N__23518\,
            I => \N__23514\
        );

    \I__2934\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23511\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__23514\,
            I => \N__23508\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__23511\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__2931\ : Odrv4
    port map (
            O => \N__23508\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__2930\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23500\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__23500\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\
        );

    \I__2928\ : InMux
    port map (
            O => \N__23497\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__2927\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23490\
        );

    \I__2926\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23487\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__23490\,
            I => \N__23484\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__23487\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__23484\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__23479\,
            I => \N__23476\
        );

    \I__2921\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23473\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__23473\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\
        );

    \I__2919\ : InMux
    port map (
            O => \N__23470\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__23467\,
            I => \N__23463\
        );

    \I__2917\ : InMux
    port map (
            O => \N__23466\,
            I => \N__23460\
        );

    \I__2916\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23457\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23454\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__23457\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__23454\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__2912\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23446\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__23446\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\
        );

    \I__2910\ : InMux
    port map (
            O => \N__23443\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__2909\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23436\
        );

    \I__2908\ : InMux
    port map (
            O => \N__23439\,
            I => \N__23433\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__23436\,
            I => \N__23430\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__23433\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__23430\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__23425\,
            I => \N__23422\
        );

    \I__2903\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23419\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__23419\,
            I => \N__23416\
        );

    \I__2901\ : Span4Mux_h
    port map (
            O => \N__23416\,
            I => \N__23413\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__23413\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\
        );

    \I__2899\ : InMux
    port map (
            O => \N__23410\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__2898\ : InMux
    port map (
            O => \N__23407\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__23404\,
            I => \N__23401\
        );

    \I__2896\ : InMux
    port map (
            O => \N__23401\,
            I => \N__23398\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__23398\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__23395\,
            I => \N__23392\
        );

    \I__2893\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23389\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__23389\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__23386\,
            I => \N__23383\
        );

    \I__2890\ : InMux
    port map (
            O => \N__23383\,
            I => \N__23380\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__23380\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__23377\,
            I => \N__23372\
        );

    \I__2887\ : InMux
    port map (
            O => \N__23376\,
            I => \N__23369\
        );

    \I__2886\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23366\
        );

    \I__2885\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23363\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__23369\,
            I => \N__23360\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__23366\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__23363\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__23360\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__2880\ : InMux
    port map (
            O => \N__23353\,
            I => \N__23350\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__23350\,
            I => \N__23346\
        );

    \I__2878\ : InMux
    port map (
            O => \N__23349\,
            I => \N__23343\
        );

    \I__2877\ : Span4Mux_h
    port map (
            O => \N__23346\,
            I => \N__23340\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__23343\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__2875\ : Odrv4
    port map (
            O => \N__23340\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__2874\ : InMux
    port map (
            O => \N__23335\,
            I => \N__23332\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__23332\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\
        );

    \I__2872\ : InMux
    port map (
            O => \N__23329\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__2871\ : InMux
    port map (
            O => \N__23326\,
            I => \N__23322\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__23325\,
            I => \N__23319\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__23322\,
            I => \N__23316\
        );

    \I__2868\ : InMux
    port map (
            O => \N__23319\,
            I => \N__23313\
        );

    \I__2867\ : Span4Mux_h
    port map (
            O => \N__23316\,
            I => \N__23310\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__23313\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__2865\ : Odrv4
    port map (
            O => \N__23310\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__2864\ : InMux
    port map (
            O => \N__23305\,
            I => \N__23302\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__23302\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\
        );

    \I__2862\ : InMux
    port map (
            O => \N__23299\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__2861\ : InMux
    port map (
            O => \N__23296\,
            I => \N__23293\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__23293\,
            I => \N__23289\
        );

    \I__2859\ : InMux
    port map (
            O => \N__23292\,
            I => \N__23286\
        );

    \I__2858\ : Span4Mux_h
    port map (
            O => \N__23289\,
            I => \N__23283\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__23286\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__2856\ : Odrv4
    port map (
            O => \N__23283\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__2855\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23275\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__23275\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\
        );

    \I__2853\ : InMux
    port map (
            O => \N__23272\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__2852\ : InMux
    port map (
            O => \N__23269\,
            I => \N__23265\
        );

    \I__2851\ : InMux
    port map (
            O => \N__23268\,
            I => \N__23262\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__23265\,
            I => \N__23257\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__23262\,
            I => \N__23257\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__23257\,
            I => \N__23254\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__23254\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__2846\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23248\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__23248\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__2844\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23242\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__23242\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__2842\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23236\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__23236\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__2840\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23230\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__23230\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__23227\,
            I => \N__23224\
        );

    \I__2837\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23221\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__23221\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__2835\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23215\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__23215\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__2833\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23209\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__23209\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__2831\ : InMux
    port map (
            O => \N__23206\,
            I => \N__23203\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__23203\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__2829\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23197\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__23197\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__2827\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23191\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__23191\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__2825\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23185\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__23185\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__2823\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23179\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__23179\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__2821\ : InMux
    port map (
            O => \N__23176\,
            I => \N__23173\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__23173\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__23170\,
            I => \N__23167\
        );

    \I__2818\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23164\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__23164\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__2816\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23158\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__23158\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__2814\ : InMux
    port map (
            O => \N__23155\,
            I => \N__23152\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__23152\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__2812\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23146\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__23146\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__23143\,
            I => \N__23140\
        );

    \I__2809\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23137\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__23137\,
            I => \N__23134\
        );

    \I__2807\ : Odrv12
    port map (
            O => \N__23134\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__2806\ : InMux
    port map (
            O => \N__23131\,
            I => \N__23128\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__23128\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__2804\ : InMux
    port map (
            O => \N__23125\,
            I => \N__23122\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__23122\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__23119\,
            I => \N__23116\
        );

    \I__2801\ : InMux
    port map (
            O => \N__23116\,
            I => \N__23113\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__23113\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17\
        );

    \I__2799\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23107\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__23107\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__23104\,
            I => \N__23101\
        );

    \I__2796\ : InMux
    port map (
            O => \N__23101\,
            I => \N__23098\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__23098\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19\
        );

    \I__2794\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23092\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__23092\,
            I => \N__23089\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__23089\,
            I => \N__23086\
        );

    \I__2791\ : Odrv4
    port map (
            O => \N__23086\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__2790\ : InMux
    port map (
            O => \N__23083\,
            I => \N__23080\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__23080\,
            I => \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__23077\,
            I => \N__23074\
        );

    \I__2787\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__23071\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9\
        );

    \I__2785\ : InMux
    port map (
            O => \N__23068\,
            I => \N__23065\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__23065\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16\
        );

    \I__2783\ : InMux
    port map (
            O => \N__23062\,
            I => \N__23059\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__23059\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__2781\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23053\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__23053\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__2779\ : InMux
    port map (
            O => \N__23050\,
            I => \N__23047\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__23047\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__23044\,
            I => \phase_controller_inst2.stoper_tr.time_passed11_cascade_\
        );

    \I__2776\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23038\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__23038\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0\
        );

    \I__2774\ : InMux
    port map (
            O => \N__23035\,
            I => \N__23030\
        );

    \I__2773\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23027\
        );

    \I__2772\ : InMux
    port map (
            O => \N__23033\,
            I => \N__23024\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__23030\,
            I => \phase_controller_inst2.stoper_tr.time_passed11\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__23027\,
            I => \phase_controller_inst2.stoper_tr.time_passed11\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__23024\,
            I => \phase_controller_inst2.stoper_tr.time_passed11\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__23017\,
            I => \N__23014\
        );

    \I__2767\ : InMux
    port map (
            O => \N__23014\,
            I => \N__23011\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__23011\,
            I => \N__23008\
        );

    \I__2765\ : Odrv4
    port map (
            O => \N__23008\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__23005\,
            I => \N__23002\
        );

    \I__2763\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22999\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__22999\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10\
        );

    \I__2761\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22993\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__22993\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11\
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__22990\,
            I => \N__22987\
        );

    \I__2758\ : InMux
    port map (
            O => \N__22987\,
            I => \N__22984\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__22984\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12\
        );

    \I__2756\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22978\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__22978\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__22975\,
            I => \N__22972\
        );

    \I__2753\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22969\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__22969\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14\
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__22966\,
            I => \N__22963\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22963\,
            I => \N__22960\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__22960\,
            I => \N__22957\
        );

    \I__2748\ : Span4Mux_h
    port map (
            O => \N__22957\,
            I => \N__22954\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__22954\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7\
        );

    \I__2746\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22948\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__22948\,
            I => \N__22945\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__22945\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3\
        );

    \I__2743\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22939\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__22939\,
            I => \N__22936\
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__22936\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2\
        );

    \I__2740\ : InMux
    port map (
            O => \N__22933\,
            I => \N__22930\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__22930\,
            I => \N__22927\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__22927\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__22924\,
            I => \N__22921\
        );

    \I__2736\ : InMux
    port map (
            O => \N__22921\,
            I => \N__22918\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__22918\,
            I => \N__22915\
        );

    \I__2734\ : Span4Mux_h
    port map (
            O => \N__22915\,
            I => \N__22912\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__22912\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6\
        );

    \I__2732\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22906\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__22906\,
            I => \N__22903\
        );

    \I__2730\ : Odrv4
    port map (
            O => \N__22903\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__22900\,
            I => \N__22897\
        );

    \I__2728\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22894\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__22894\,
            I => \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__22891\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\
        );

    \I__2725\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22885\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__22885\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2723\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22879\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__22879\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__22876\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__2720\ : InMux
    port map (
            O => \N__22873\,
            I => \N__22870\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__22870\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2718\ : InMux
    port map (
            O => \N__22867\,
            I => \N__22864\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__22864\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2716\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22858\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__22858\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2714\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22852\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__22852\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\
        );

    \I__2712\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22846\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__22846\,
            I => \N__22843\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__22843\,
            I => il_max_comp1_c
        );

    \I__2709\ : InMux
    port map (
            O => \N__22840\,
            I => \N__22837\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__22837\,
            I => \il_max_comp1_D1\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__22834\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\
        );

    \I__2706\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22828\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__22828\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__22825\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__22822\,
            I => \N__22817\
        );

    \I__2702\ : InMux
    port map (
            O => \N__22821\,
            I => \N__22807\
        );

    \I__2701\ : InMux
    port map (
            O => \N__22820\,
            I => \N__22807\
        );

    \I__2700\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22800\
        );

    \I__2699\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22800\
        );

    \I__2698\ : InMux
    port map (
            O => \N__22815\,
            I => \N__22800\
        );

    \I__2697\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22797\
        );

    \I__2696\ : InMux
    port map (
            O => \N__22813\,
            I => \N__22792\
        );

    \I__2695\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22792\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__22807\,
            I => \N__22789\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__22800\,
            I => \N__22786\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__22797\,
            I => \N__22781\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__22792\,
            I => \N__22781\
        );

    \I__2690\ : Span4Mux_h
    port map (
            O => \N__22789\,
            I => \N__22778\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__22786\,
            I => \N__22775\
        );

    \I__2688\ : Span4Mux_h
    port map (
            O => \N__22781\,
            I => \N__22772\
        );

    \I__2687\ : Span4Mux_v
    port map (
            O => \N__22778\,
            I => \N__22769\
        );

    \I__2686\ : Span4Mux_h
    port map (
            O => \N__22775\,
            I => \N__22766\
        );

    \I__2685\ : Span4Mux_h
    port map (
            O => \N__22772\,
            I => \N__22763\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__22769\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2683\ : Odrv4
    port map (
            O => \N__22766\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__22763\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2681\ : InMux
    port map (
            O => \N__22756\,
            I => \N__22753\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__22753\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__22750\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\
        );

    \I__2678\ : InMux
    port map (
            O => \N__22747\,
            I => \N__22735\
        );

    \I__2677\ : InMux
    port map (
            O => \N__22746\,
            I => \N__22735\
        );

    \I__2676\ : InMux
    port map (
            O => \N__22745\,
            I => \N__22735\
        );

    \I__2675\ : InMux
    port map (
            O => \N__22744\,
            I => \N__22730\
        );

    \I__2674\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22730\
        );

    \I__2673\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22727\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22723\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22718\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__22727\,
            I => \N__22718\
        );

    \I__2669\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22715\
        );

    \I__2668\ : Span4Mux_h
    port map (
            O => \N__22723\,
            I => \N__22712\
        );

    \I__2667\ : Sp12to4
    port map (
            O => \N__22718\,
            I => \N__22707\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__22715\,
            I => \N__22707\
        );

    \I__2665\ : Span4Mux_h
    port map (
            O => \N__22712\,
            I => \N__22704\
        );

    \I__2664\ : Span12Mux_s8_v
    port map (
            O => \N__22707\,
            I => \N__22701\
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__22704\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2662\ : Odrv12
    port map (
            O => \N__22701\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2661\ : InMux
    port map (
            O => \N__22696\,
            I => \N__22693\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__22693\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2659\ : InMux
    port map (
            O => \N__22690\,
            I => \N__22687\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__22687\,
            I => \N__22682\
        );

    \I__2657\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22679\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__22685\,
            I => \N__22676\
        );

    \I__2655\ : Span12Mux_v
    port map (
            O => \N__22682\,
            I => \N__22670\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__22679\,
            I => \N__22670\
        );

    \I__2653\ : InMux
    port map (
            O => \N__22676\,
            I => \N__22667\
        );

    \I__2652\ : InMux
    port map (
            O => \N__22675\,
            I => \N__22664\
        );

    \I__2651\ : Odrv12
    port map (
            O => \N__22670\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__22667\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22664\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__2648\ : IoInMux
    port map (
            O => \N__22657\,
            I => \N__22654\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__22654\,
            I => \N__22651\
        );

    \I__2646\ : Span12Mux_s7_v
    port map (
            O => \N__22651\,
            I => \N__22648\
        );

    \I__2645\ : Odrv12
    port map (
            O => \N__22648\,
            I => s4_phy_c
        );

    \I__2644\ : InMux
    port map (
            O => \N__22645\,
            I => \N__22642\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__22642\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\
        );

    \I__2642\ : InMux
    port map (
            O => \N__22639\,
            I => \bfn_7_17_0_\
        );

    \I__2641\ : InMux
    port map (
            O => \N__22636\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__2640\ : InMux
    port map (
            O => \N__22633\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__2639\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22626\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__22629\,
            I => \N__22622\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__22626\,
            I => \N__22619\
        );

    \I__2636\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22616\
        );

    \I__2635\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22613\
        );

    \I__2634\ : Span4Mux_h
    port map (
            O => \N__22619\,
            I => \N__22610\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__22616\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__22613\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__22610\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__22603\,
            I => \N__22600\
        );

    \I__2629\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22597\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__22597\,
            I => \N__22594\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__22594\,
            I => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__2626\ : InMux
    port map (
            O => \N__22591\,
            I => \N__22588\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__22588\,
            I => \N__22584\
        );

    \I__2624\ : InMux
    port map (
            O => \N__22587\,
            I => \N__22581\
        );

    \I__2623\ : Span4Mux_h
    port map (
            O => \N__22584\,
            I => \N__22575\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__22581\,
            I => \N__22575\
        );

    \I__2621\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22572\
        );

    \I__2620\ : Span4Mux_v
    port map (
            O => \N__22575\,
            I => \N__22569\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__22572\,
            I => \N__22566\
        );

    \I__2618\ : Span4Mux_v
    port map (
            O => \N__22569\,
            I => \N__22563\
        );

    \I__2617\ : Odrv12
    port map (
            O => \N__22566\,
            I => \il_min_comp1_D2\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__22563\,
            I => \il_min_comp1_D2\
        );

    \I__2615\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22553\
        );

    \I__2614\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22550\
        );

    \I__2613\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22547\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22544\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__22550\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__22547\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__2609\ : Odrv4
    port map (
            O => \N__22544\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__2608\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22533\
        );

    \I__2607\ : InMux
    port map (
            O => \N__22536\,
            I => \N__22530\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__22533\,
            I => \N__22527\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__22530\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__22527\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__2603\ : InMux
    port map (
            O => \N__22522\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__2602\ : InMux
    port map (
            O => \N__22519\,
            I => \bfn_7_16_0_\
        );

    \I__2601\ : InMux
    port map (
            O => \N__22516\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__2600\ : InMux
    port map (
            O => \N__22513\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__2599\ : InMux
    port map (
            O => \N__22510\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__2598\ : InMux
    port map (
            O => \N__22507\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__2597\ : InMux
    port map (
            O => \N__22504\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__2596\ : InMux
    port map (
            O => \N__22501\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__2595\ : InMux
    port map (
            O => \N__22498\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__22495\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__22492\,
            I => \N__22488\
        );

    \I__2592\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22485\
        );

    \I__2591\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22482\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__22485\,
            I => \N__22479\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__22482\,
            I => \N__22476\
        );

    \I__2588\ : Odrv4
    port map (
            O => \N__22479\,
            I => state_ns_i_a3_1
        );

    \I__2587\ : Odrv12
    port map (
            O => \N__22476\,
            I => state_ns_i_a3_1
        );

    \I__2586\ : InMux
    port map (
            O => \N__22471\,
            I => \N__22466\
        );

    \I__2585\ : InMux
    port map (
            O => \N__22470\,
            I => \N__22463\
        );

    \I__2584\ : InMux
    port map (
            O => \N__22469\,
            I => \N__22460\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__22466\,
            I => \N__22453\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__22463\,
            I => \N__22453\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__22460\,
            I => \N__22453\
        );

    \I__2580\ : Odrv12
    port map (
            O => \N__22453\,
            I => \il_min_comp2_D2\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__22450\,
            I => \N__22447\
        );

    \I__2578\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22440\
        );

    \I__2577\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22440\
        );

    \I__2576\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22437\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__22440\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__22437\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__2573\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22426\
        );

    \I__2572\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22426\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__22426\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__2570\ : InMux
    port map (
            O => \N__22423\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__2569\ : InMux
    port map (
            O => \N__22420\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__2568\ : InMux
    port map (
            O => \N__22417\,
            I => \N__22414\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__22414\,
            I => \N__22411\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__22411\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4\
        );

    \I__2565\ : InMux
    port map (
            O => \N__22408\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__2564\ : InMux
    port map (
            O => \N__22405\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__2563\ : InMux
    port map (
            O => \N__22402\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__2562\ : InMux
    port map (
            O => \N__22399\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__2561\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22393\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22390\
        );

    \I__2559\ : Span4Mux_h
    port map (
            O => \N__22390\,
            I => \N__22387\
        );

    \I__2558\ : Span4Mux_v
    port map (
            O => \N__22387\,
            I => \N__22384\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__22384\,
            I => il_max_comp2_c
        );

    \I__2556\ : InMux
    port map (
            O => \N__22381\,
            I => \N__22378\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__22378\,
            I => \N__22375\
        );

    \I__2554\ : Odrv4
    port map (
            O => \N__22375\,
            I => \il_max_comp2_D1\
        );

    \I__2553\ : IoInMux
    port map (
            O => \N__22372\,
            I => \N__22369\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__22369\,
            I => \N__22366\
        );

    \I__2551\ : IoSpan4Mux
    port map (
            O => \N__22366\,
            I => \N__22363\
        );

    \I__2550\ : Span4Mux_s1_v
    port map (
            O => \N__22363\,
            I => \N__22360\
        );

    \I__2549\ : Sp12to4
    port map (
            O => \N__22360\,
            I => \N__22357\
        );

    \I__2548\ : Span12Mux_s9_v
    port map (
            O => \N__22357\,
            I => \N__22354\
        );

    \I__2547\ : Odrv12
    port map (
            O => \N__22354\,
            I => \delay_measurement_inst.delay_hc_timer.N_302_i\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__22351\,
            I => \N__22348\
        );

    \I__2545\ : InMux
    port map (
            O => \N__22348\,
            I => \N__22345\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__22345\,
            I => \phase_controller_inst2.start_timer_tr_0_sqmuxa\
        );

    \I__2543\ : InMux
    port map (
            O => \N__22342\,
            I => \N__22339\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__22339\,
            I => \N__22336\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__22336\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__2540\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22329\
        );

    \I__2539\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22326\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__22329\,
            I => \N__22321\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__22326\,
            I => \N__22321\
        );

    \I__2536\ : Span4Mux_s3_v
    port map (
            O => \N__22321\,
            I => \N__22318\
        );

    \I__2535\ : Span4Mux_h
    port map (
            O => \N__22318\,
            I => \N__22313\
        );

    \I__2534\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22310\
        );

    \I__2533\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22307\
        );

    \I__2532\ : Sp12to4
    port map (
            O => \N__22313\,
            I => \N__22304\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__22310\,
            I => \N__22299\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22299\
        );

    \I__2529\ : Span12Mux_v
    port map (
            O => \N__22304\,
            I => \N__22294\
        );

    \I__2528\ : Sp12to4
    port map (
            O => \N__22299\,
            I => \N__22294\
        );

    \I__2527\ : Span12Mux_v
    port map (
            O => \N__22294\,
            I => \N__22291\
        );

    \I__2526\ : Span12Mux_h
    port map (
            O => \N__22291\,
            I => \N__22288\
        );

    \I__2525\ : Odrv12
    port map (
            O => \N__22288\,
            I => start_stop_c
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__22285\,
            I => \N__22282\
        );

    \I__2523\ : InMux
    port map (
            O => \N__22282\,
            I => \N__22279\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__22279\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__2521\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22273\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__22273\,
            I => \N__22269\
        );

    \I__2519\ : InMux
    port map (
            O => \N__22272\,
            I => \N__22266\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__22269\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__22266\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__2516\ : InMux
    port map (
            O => \N__22261\,
            I => \N__22254\
        );

    \I__2515\ : InMux
    port map (
            O => \N__22260\,
            I => \N__22254\
        );

    \I__2514\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22251\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__22254\,
            I => \N__22248\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__22251\,
            I => \N__22245\
        );

    \I__2511\ : Span4Mux_h
    port map (
            O => \N__22248\,
            I => \N__22242\
        );

    \I__2510\ : Span4Mux_h
    port map (
            O => \N__22245\,
            I => \N__22239\
        );

    \I__2509\ : Sp12to4
    port map (
            O => \N__22242\,
            I => \N__22236\
        );

    \I__2508\ : Span4Mux_v
    port map (
            O => \N__22239\,
            I => \N__22233\
        );

    \I__2507\ : Span12Mux_v
    port map (
            O => \N__22236\,
            I => \N__22230\
        );

    \I__2506\ : Span4Mux_v
    port map (
            O => \N__22233\,
            I => \N__22227\
        );

    \I__2505\ : Odrv12
    port map (
            O => \N__22230\,
            I => \il_max_comp1_D2\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__22227\,
            I => \il_max_comp1_D2\
        );

    \I__2503\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22219\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__22219\,
            I => \N__22216\
        );

    \I__2501\ : Odrv12
    port map (
            O => \N__22216\,
            I => il_min_comp2_c
        );

    \I__2500\ : InMux
    port map (
            O => \N__22213\,
            I => \N__22210\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__22210\,
            I => \il_min_comp2_D1\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__22207\,
            I => \N__22204\
        );

    \I__2497\ : InMux
    port map (
            O => \N__22204\,
            I => \N__22201\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__22201\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__2495\ : InMux
    port map (
            O => \N__22198\,
            I => \N__22193\
        );

    \I__2494\ : InMux
    port map (
            O => \N__22197\,
            I => \N__22190\
        );

    \I__2493\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22187\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__22193\,
            I => \N__22182\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__22190\,
            I => \N__22182\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__22187\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__22182\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2488\ : InMux
    port map (
            O => \N__22177\,
            I => \N__22174\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__22174\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2486\ : InMux
    port map (
            O => \N__22171\,
            I => \N__22166\
        );

    \I__2485\ : InMux
    port map (
            O => \N__22170\,
            I => \N__22163\
        );

    \I__2484\ : InMux
    port map (
            O => \N__22169\,
            I => \N__22160\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__22166\,
            I => \N__22155\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__22163\,
            I => \N__22155\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__22160\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__22155\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2479\ : CascadeMux
    port map (
            O => \N__22150\,
            I => \N__22147\
        );

    \I__2478\ : InMux
    port map (
            O => \N__22147\,
            I => \N__22144\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__22144\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__2476\ : InMux
    port map (
            O => \N__22141\,
            I => \N__22138\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__22138\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__2473\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22129\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__22129\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__2471\ : InMux
    port map (
            O => \N__22126\,
            I => \N__22121\
        );

    \I__2470\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22118\
        );

    \I__2469\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22115\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__22121\,
            I => \N__22112\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__22118\,
            I => \N__22109\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__22115\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__22112\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__22109\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2463\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22099\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__22099\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__22096\,
            I => \N__22093\
        );

    \I__2460\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22090\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__22090\,
            I => \N__22087\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__22087\,
            I => \N__22084\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__22084\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__2456\ : InMux
    port map (
            O => \N__22081\,
            I => \N__22076\
        );

    \I__2455\ : InMux
    port map (
            O => \N__22080\,
            I => \N__22073\
        );

    \I__2454\ : InMux
    port map (
            O => \N__22079\,
            I => \N__22070\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__22076\,
            I => \N__22067\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22064\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__22070\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2450\ : Odrv12
    port map (
            O => \N__22067\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__22064\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2448\ : InMux
    port map (
            O => \N__22057\,
            I => \N__22054\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__22054\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__22051\,
            I => \N__22048\
        );

    \I__2445\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22045\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__22045\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__2443\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22037\
        );

    \I__2442\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22034\
        );

    \I__2441\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22031\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__22037\,
            I => \N__22028\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__22034\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__22031\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2437\ : Odrv12
    port map (
            O => \N__22028\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2436\ : InMux
    port map (
            O => \N__22021\,
            I => \N__22018\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__22018\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2434\ : InMux
    port map (
            O => \N__22015\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2433\ : IoInMux
    port map (
            O => \N__22012\,
            I => \N__22009\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__2431\ : Span4Mux_s1_v
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__2430\ : Span4Mux_h
    port map (
            O => \N__22003\,
            I => \N__22000\
        );

    \I__2429\ : Sp12to4
    port map (
            O => \N__22000\,
            I => \N__21997\
        );

    \I__2428\ : Span12Mux_h
    port map (
            O => \N__21997\,
            I => \N__21994\
        );

    \I__2427\ : Odrv12
    port map (
            O => \N__21994\,
            I => pwm_output_c
        );

    \I__2426\ : CascadeMux
    port map (
            O => \N__21991\,
            I => \pwm_generator_inst.un1_counterlto9_2_cascade_\
        );

    \I__2425\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21970\
        );

    \I__2424\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21970\
        );

    \I__2423\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21970\
        );

    \I__2422\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21970\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21984\,
            I => \N__21961\
        );

    \I__2420\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21961\
        );

    \I__2419\ : InMux
    port map (
            O => \N__21982\,
            I => \N__21961\
        );

    \I__2418\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21961\
        );

    \I__2417\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21956\
        );

    \I__2416\ : InMux
    port map (
            O => \N__21979\,
            I => \N__21956\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__21970\,
            I => \N__21951\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__21961\,
            I => \N__21951\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__21956\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2412\ : Odrv4
    port map (
            O => \N__21951\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__21946\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__2410\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21940\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__21940\,
            I => \pwm_generator_inst.un1_counterlt9\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__21937\,
            I => \N__21934\
        );

    \I__2407\ : InMux
    port map (
            O => \N__21934\,
            I => \N__21931\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__21931\,
            I => \N__21928\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__21928\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21920\
        );

    \I__2403\ : InMux
    port map (
            O => \N__21924\,
            I => \N__21917\
        );

    \I__2402\ : InMux
    port map (
            O => \N__21923\,
            I => \N__21914\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__21920\,
            I => \N__21911\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__21917\,
            I => \N__21908\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__21914\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2398\ : Odrv12
    port map (
            O => \N__21911\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2397\ : Odrv4
    port map (
            O => \N__21908\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2396\ : InMux
    port map (
            O => \N__21901\,
            I => \N__21898\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__21898\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__21895\,
            I => \N__21892\
        );

    \I__2393\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21889\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__21889\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__2391\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21881\
        );

    \I__2390\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21878\
        );

    \I__2389\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21875\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__21881\,
            I => \N__21872\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__21878\,
            I => \N__21869\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__21875\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2385\ : Odrv12
    port map (
            O => \N__21872\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__21869\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2383\ : InMux
    port map (
            O => \N__21862\,
            I => \N__21859\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__21859\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__21856\,
            I => \N__21853\
        );

    \I__2380\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21850\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__21850\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__2378\ : InMux
    port map (
            O => \N__21847\,
            I => \N__21842\
        );

    \I__2377\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21839\
        );

    \I__2376\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21836\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__21842\,
            I => \N__21831\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__21839\,
            I => \N__21831\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__21836\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2372\ : Odrv4
    port map (
            O => \N__21831\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2371\ : InMux
    port map (
            O => \N__21826\,
            I => \N__21823\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__21823\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__21820\,
            I => \N__21817\
        );

    \I__2368\ : InMux
    port map (
            O => \N__21817\,
            I => \N__21814\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__21814\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__2366\ : InMux
    port map (
            O => \N__21811\,
            I => \N__21806\
        );

    \I__2365\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21803\
        );

    \I__2364\ : InMux
    port map (
            O => \N__21809\,
            I => \N__21800\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__21806\,
            I => \N__21795\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__21803\,
            I => \N__21795\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__21800\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2360\ : Odrv4
    port map (
            O => \N__21795\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2359\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21787\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__21787\,
            I => \N__21784\
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__21784\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__21781\,
            I => \N__21778\
        );

    \I__2355\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21775\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__21775\,
            I => \N__21772\
        );

    \I__2353\ : Span4Mux_h
    port map (
            O => \N__21772\,
            I => \N__21769\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__21769\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__2351\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21761\
        );

    \I__2350\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21758\
        );

    \I__2349\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21755\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__21761\,
            I => \N__21750\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21750\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__21755\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__21750\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2344\ : InMux
    port map (
            O => \N__21745\,
            I => \N__21742\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__21742\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2342\ : InMux
    port map (
            O => \N__21739\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__2341\ : InMux
    port map (
            O => \N__21736\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__2340\ : InMux
    port map (
            O => \N__21733\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__2339\ : InMux
    port map (
            O => \N__21730\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21727\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__2337\ : InMux
    port map (
            O => \N__21724\,
            I => \bfn_5_9_0_\
        );

    \I__2336\ : InMux
    port map (
            O => \N__21721\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__2335\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21715\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__21715\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__2333\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21709\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__21709\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__2331\ : InMux
    port map (
            O => \N__21706\,
            I => \N__21703\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__21703\,
            I => \N__21700\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__21700\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__2328\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21694\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__21694\,
            I => \N__21691\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__21691\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__2325\ : InMux
    port map (
            O => \N__21688\,
            I => \N__21685\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__21685\,
            I => \N__21682\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__21682\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__2322\ : InMux
    port map (
            O => \N__21679\,
            I => \N__21676\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__21676\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__2320\ : InMux
    port map (
            O => \N__21673\,
            I => \bfn_5_8_0_\
        );

    \I__2319\ : InMux
    port map (
            O => \N__21670\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__2318\ : InMux
    port map (
            O => \N__21667\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__2317\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21661\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__21661\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__2315\ : InMux
    port map (
            O => \N__21658\,
            I => \N__21655\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__21655\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__2313\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21649\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__21649\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__2311\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__21643\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__2309\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__21637\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__2307\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21631\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__21631\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__21628\,
            I => \N__21621\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__21627\,
            I => \N__21617\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__21626\,
            I => \N__21614\
        );

    \I__2302\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21589\
        );

    \I__2301\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21589\
        );

    \I__2300\ : InMux
    port map (
            O => \N__21621\,
            I => \N__21586\
        );

    \I__2299\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21583\
        );

    \I__2298\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21578\
        );

    \I__2297\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21578\
        );

    \I__2296\ : InMux
    port map (
            O => \N__21613\,
            I => \N__21569\
        );

    \I__2295\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21569\
        );

    \I__2294\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21569\
        );

    \I__2293\ : InMux
    port map (
            O => \N__21610\,
            I => \N__21569\
        );

    \I__2292\ : InMux
    port map (
            O => \N__21609\,
            I => \N__21551\
        );

    \I__2291\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21551\
        );

    \I__2290\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21551\
        );

    \I__2289\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21551\
        );

    \I__2288\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21551\
        );

    \I__2287\ : InMux
    port map (
            O => \N__21604\,
            I => \N__21551\
        );

    \I__2286\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21551\
        );

    \I__2285\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21551\
        );

    \I__2284\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21548\
        );

    \I__2283\ : InMux
    port map (
            O => \N__21600\,
            I => \N__21533\
        );

    \I__2282\ : InMux
    port map (
            O => \N__21599\,
            I => \N__21533\
        );

    \I__2281\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21533\
        );

    \I__2280\ : InMux
    port map (
            O => \N__21597\,
            I => \N__21533\
        );

    \I__2279\ : InMux
    port map (
            O => \N__21596\,
            I => \N__21533\
        );

    \I__2278\ : InMux
    port map (
            O => \N__21595\,
            I => \N__21533\
        );

    \I__2277\ : InMux
    port map (
            O => \N__21594\,
            I => \N__21533\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__21589\,
            I => \N__21530\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__21586\,
            I => \N__21521\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__21583\,
            I => \N__21521\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__21578\,
            I => \N__21521\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__21569\,
            I => \N__21521\
        );

    \I__2271\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21518\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__21551\,
            I => \N__21515\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__21548\,
            I => \N__21510\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__21533\,
            I => \N__21510\
        );

    \I__2267\ : Span4Mux_v
    port map (
            O => \N__21530\,
            I => \N__21500\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__21521\,
            I => \N__21500\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__21518\,
            I => \N__21497\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__21515\,
            I => \N__21492\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__21510\,
            I => \N__21492\
        );

    \I__2262\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21487\
        );

    \I__2261\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21487\
        );

    \I__2260\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21480\
        );

    \I__2259\ : InMux
    port map (
            O => \N__21506\,
            I => \N__21480\
        );

    \I__2258\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21480\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__21500\,
            I => \N_19_1\
        );

    \I__2256\ : Odrv12
    port map (
            O => \N__21497\,
            I => \N_19_1\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__21492\,
            I => \N_19_1\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__21487\,
            I => \N_19_1\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__21480\,
            I => \N_19_1\
        );

    \I__2252\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21448\
        );

    \I__2251\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21448\
        );

    \I__2250\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21448\
        );

    \I__2249\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21448\
        );

    \I__2248\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21448\
        );

    \I__2247\ : InMux
    port map (
            O => \N__21464\,
            I => \N__21448\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__21463\,
            I => \N__21445\
        );

    \I__2245\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21439\
        );

    \I__2244\ : InMux
    port map (
            O => \N__21461\,
            I => \N__21439\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__21448\,
            I => \N__21436\
        );

    \I__2242\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21431\
        );

    \I__2241\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21431\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__21439\,
            I => \N__21428\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__21436\,
            I => \N__21423\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__21431\,
            I => \N__21423\
        );

    \I__2237\ : Odrv12
    port map (
            O => \N__21428\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2236\ : Odrv4
    port map (
            O => \N__21423\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__21418\,
            I => \N__21410\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__21417\,
            I => \N__21407\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__21416\,
            I => \N__21402\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__21415\,
            I => \N__21399\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__21414\,
            I => \N__21396\
        );

    \I__2230\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21389\
        );

    \I__2229\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21389\
        );

    \I__2228\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21376\
        );

    \I__2227\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21376\
        );

    \I__2226\ : InMux
    port map (
            O => \N__21405\,
            I => \N__21376\
        );

    \I__2225\ : InMux
    port map (
            O => \N__21402\,
            I => \N__21376\
        );

    \I__2224\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21376\
        );

    \I__2223\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21376\
        );

    \I__2222\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21371\
        );

    \I__2221\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21371\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__21389\,
            I => \N__21368\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__21376\,
            I => \N__21363\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__21371\,
            I => \N__21363\
        );

    \I__2217\ : Span4Mux_v
    port map (
            O => \N__21368\,
            I => \N__21360\
        );

    \I__2216\ : Span4Mux_v
    port map (
            O => \N__21363\,
            I => \N__21357\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__21360\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__21357\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2213\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21349\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__21349\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__2211\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21343\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__21343\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__2209\ : InMux
    port map (
            O => \N__21340\,
            I => \N__21337\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__21337\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__2207\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21331\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__21331\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__2205\ : InMux
    port map (
            O => \N__21328\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__21325\,
            I => \N__21322\
        );

    \I__2203\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21319\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__21319\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__2201\ : InMux
    port map (
            O => \N__21316\,
            I => \bfn_3_9_0_\
        );

    \I__2200\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21310\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__21310\,
            I => \N__21307\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__21307\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__21304\,
            I => \N__21299\
        );

    \I__2196\ : InMux
    port map (
            O => \N__21303\,
            I => \N__21287\
        );

    \I__2195\ : InMux
    port map (
            O => \N__21302\,
            I => \N__21284\
        );

    \I__2194\ : InMux
    port map (
            O => \N__21299\,
            I => \N__21281\
        );

    \I__2193\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21272\
        );

    \I__2192\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21272\
        );

    \I__2191\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21272\
        );

    \I__2190\ : InMux
    port map (
            O => \N__21295\,
            I => \N__21272\
        );

    \I__2189\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21263\
        );

    \I__2188\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21263\
        );

    \I__2187\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21263\
        );

    \I__2186\ : InMux
    port map (
            O => \N__21291\,
            I => \N__21263\
        );

    \I__2185\ : InMux
    port map (
            O => \N__21290\,
            I => \N__21260\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__21287\,
            I => \N__21253\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__21284\,
            I => \N__21253\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__21281\,
            I => \N__21253\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__21272\,
            I => \N__21246\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__21263\,
            I => \N__21246\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__21260\,
            I => \N__21246\
        );

    \I__2178\ : Span4Mux_v
    port map (
            O => \N__21253\,
            I => \N__21243\
        );

    \I__2177\ : Span4Mux_v
    port map (
            O => \N__21246\,
            I => \N__21240\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__21243\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__21240\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__21235\,
            I => \N__21232\
        );

    \I__2173\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21229\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__21229\,
            I => \N__21226\
        );

    \I__2171\ : Span4Mux_h
    port map (
            O => \N__21226\,
            I => \N__21223\
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__21223\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__2169\ : InMux
    port map (
            O => \N__21220\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__21217\,
            I => \N__21214\
        );

    \I__2167\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21211\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__21211\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__2165\ : InMux
    port map (
            O => \N__21208\,
            I => \N__21205\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__21205\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__2163\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21199\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__21199\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__2161\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21193\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__21193\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__2159\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21187\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__21187\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__21184\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__2156\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21174\
        );

    \I__2155\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21174\
        );

    \I__2154\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21171\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__21174\,
            I => \N__21168\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__21171\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__21168\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2150\ : InMux
    port map (
            O => \N__21163\,
            I => \N__21160\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__21160\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__2148\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21154\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__21154\,
            I => \N__21151\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__21151\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__2145\ : InMux
    port map (
            O => \N__21148\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__2144\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21142\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__21142\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__2142\ : InMux
    port map (
            O => \N__21139\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__2141\ : InMux
    port map (
            O => \N__21136\,
            I => \N__21133\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__21133\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__2139\ : InMux
    port map (
            O => \N__21130\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__2138\ : InMux
    port map (
            O => \N__21127\,
            I => \N__21124\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__21124\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__2136\ : InMux
    port map (
            O => \N__21121\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__2135\ : InMux
    port map (
            O => \N__21118\,
            I => \N__21115\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__21115\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__2133\ : InMux
    port map (
            O => \N__21112\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__2132\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21106\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__21106\,
            I => \N__21103\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__21103\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__2129\ : InMux
    port map (
            O => \N__21100\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__2128\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21094\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__21094\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__2126\ : InMux
    port map (
            O => \N__21091\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__2125\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21085\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__21085\,
            I => \N__21082\
        );

    \I__2123\ : Span4Mux_v
    port map (
            O => \N__21082\,
            I => \N__21079\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__21079\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__2121\ : InMux
    port map (
            O => \N__21076\,
            I => \N__21073\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__21073\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__2119\ : InMux
    port map (
            O => \N__21070\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__21067\,
            I => \N__21064\
        );

    \I__2117\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21061\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__21061\,
            I => \N__21058\
        );

    \I__2115\ : Span4Mux_h
    port map (
            O => \N__21058\,
            I => \N__21055\
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__21055\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__2113\ : InMux
    port map (
            O => \N__21052\,
            I => \N__21049\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__21049\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__2111\ : InMux
    port map (
            O => \N__21046\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__2110\ : InMux
    port map (
            O => \N__21043\,
            I => \N__21040\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__21040\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__2108\ : InMux
    port map (
            O => \N__21037\,
            I => \N__21030\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__21036\,
            I => \N__21027\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__21035\,
            I => \N__21023\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__21034\,
            I => \N__21019\
        );

    \I__2104\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21015\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__21030\,
            I => \N__21012\
        );

    \I__2102\ : InMux
    port map (
            O => \N__21027\,
            I => \N__20999\
        );

    \I__2101\ : InMux
    port map (
            O => \N__21026\,
            I => \N__20999\
        );

    \I__2100\ : InMux
    port map (
            O => \N__21023\,
            I => \N__20999\
        );

    \I__2099\ : InMux
    port map (
            O => \N__21022\,
            I => \N__20999\
        );

    \I__2098\ : InMux
    port map (
            O => \N__21019\,
            I => \N__20999\
        );

    \I__2097\ : InMux
    port map (
            O => \N__21018\,
            I => \N__20999\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__21015\,
            I => \N__20992\
        );

    \I__2095\ : Span4Mux_v
    port map (
            O => \N__21012\,
            I => \N__20992\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20992\
        );

    \I__2093\ : Span4Mux_v
    port map (
            O => \N__20992\,
            I => \N__20989\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__20989\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__2091\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20983\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__20983\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20980\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20977\,
            I => \N__20974\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__20974\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__20971\,
            I => \N__20968\
        );

    \I__2085\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20965\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__20965\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20962\,
            I => \bfn_2_13_0_\
        );

    \I__2082\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20956\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__20956\,
            I => \N__20953\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__20953\,
            I => \rgb_drv_RNOZ0\
        );

    \I__2079\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20947\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__20947\,
            I => \N__20944\
        );

    \I__2077\ : Odrv4
    port map (
            O => \N__20944\,
            I => \current_shift_inst.PI_CTRL.N_162\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20938\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__20938\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__2074\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20930\
        );

    \I__2073\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20927\
        );

    \I__2072\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20924\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__20930\,
            I => \N__20919\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__20927\,
            I => \N__20919\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__20924\,
            I => \N__20916\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__20919\,
            I => pwm_duty_input_3
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__20916\,
            I => pwm_duty_input_3
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__20911\,
            I => \N__20908\
        );

    \I__2065\ : InMux
    port map (
            O => \N__20908\,
            I => \N__20905\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__20905\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__2063\ : InMux
    port map (
            O => \N__20902\,
            I => \N__20897\
        );

    \I__2062\ : InMux
    port map (
            O => \N__20901\,
            I => \N__20894\
        );

    \I__2061\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20891\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__20897\,
            I => \N__20888\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__20894\,
            I => \N__20883\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__20891\,
            I => \N__20883\
        );

    \I__2057\ : Span4Mux_s1_h
    port map (
            O => \N__20888\,
            I => \N__20880\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__20883\,
            I => pwm_duty_input_4
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__20880\,
            I => pwm_duty_input_4
        );

    \I__2054\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20872\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__20872\,
            I => \N__20869\
        );

    \I__2052\ : Span4Mux_v
    port map (
            O => \N__20869\,
            I => \N__20866\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__20866\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__20863\,
            I => \N__20860\
        );

    \I__2049\ : InMux
    port map (
            O => \N__20860\,
            I => \N__20857\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__20857\,
            I => \N__20854\
        );

    \I__2047\ : Span4Mux_v
    port map (
            O => \N__20854\,
            I => \N__20851\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__20851\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__2045\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20845\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__20845\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__2043\ : InMux
    port map (
            O => \N__20842\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__2042\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20836\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__20836\,
            I => \N__20833\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__20833\,
            I => \N__20830\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__20830\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__20827\,
            I => \N__20824\
        );

    \I__2037\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20821\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__20821\,
            I => \N__20818\
        );

    \I__2035\ : Span4Mux_h
    port map (
            O => \N__20818\,
            I => \N__20815\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__20815\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__2033\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20809\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__20809\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__2031\ : InMux
    port map (
            O => \N__20806\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__2030\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20800\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__20800\,
            I => \N__20797\
        );

    \I__2028\ : Span4Mux_v
    port map (
            O => \N__20797\,
            I => \N__20794\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__20794\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__20791\,
            I => \N__20788\
        );

    \I__2025\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20785\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__20785\,
            I => \N__20782\
        );

    \I__2023\ : Span4Mux_h
    port map (
            O => \N__20782\,
            I => \N__20779\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__20779\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__2021\ : InMux
    port map (
            O => \N__20776\,
            I => \N__20773\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__20773\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__2019\ : InMux
    port map (
            O => \N__20770\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__2018\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20764\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20761\
        );

    \I__2016\ : Span4Mux_h
    port map (
            O => \N__20761\,
            I => \N__20758\
        );

    \I__2015\ : Span4Mux_v
    port map (
            O => \N__20758\,
            I => \N__20755\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__20755\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__20752\,
            I => \N__20749\
        );

    \I__2012\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20746\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__20746\,
            I => \N__20743\
        );

    \I__2010\ : Span4Mux_h
    port map (
            O => \N__20743\,
            I => \N__20740\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__20740\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__2008\ : InMux
    port map (
            O => \N__20737\,
            I => \N__20734\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__20734\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__2006\ : InMux
    port map (
            O => \N__20731\,
            I => \bfn_2_12_0_\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20725\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__20725\,
            I => \N__20722\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__20722\,
            I => \N__20719\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__20719\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__20716\,
            I => \N__20713\
        );

    \I__2000\ : InMux
    port map (
            O => \N__20713\,
            I => \N__20710\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__20710\,
            I => \N__20707\
        );

    \I__1998\ : Span4Mux_h
    port map (
            O => \N__20707\,
            I => \N__20704\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__20704\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1996\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20698\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__20698\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__1994\ : InMux
    port map (
            O => \N__20695\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__20692\,
            I => \N__20689\
        );

    \I__1992\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20686\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__20686\,
            I => \N__20683\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__20683\,
            I => \N__20680\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__20680\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1988\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20674\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__20674\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20671\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1985\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20665\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__20665\,
            I => \N__20662\
        );

    \I__1983\ : Span4Mux_h
    port map (
            O => \N__20662\,
            I => \N__20659\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__20659\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1981\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20653\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__20653\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__1979\ : InMux
    port map (
            O => \N__20650\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__1977\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20641\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__20641\,
            I => \N__20638\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__20638\,
            I => \N__20635\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__20635\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1973\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20628\
        );

    \I__1972\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20625\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__20628\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__20625\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1969\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20614\
        );

    \I__1968\ : InMux
    port map (
            O => \N__20619\,
            I => \N__20614\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__20614\,
            I => \N__20611\
        );

    \I__1966\ : Span4Mux_h
    port map (
            O => \N__20611\,
            I => \N__20608\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__20608\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1964\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20602\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__20602\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__20599\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\
        );

    \I__1961\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20593\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__20593\,
            I => \N__20589\
        );

    \I__1959\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20586\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__20589\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__20586\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__1956\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20577\
        );

    \I__1955\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20573\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20570\
        );

    \I__1953\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20567\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__20573\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__20570\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__20567\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__1949\ : InMux
    port map (
            O => \N__20560\,
            I => \N__20557\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__20557\,
            I => \N__20554\
        );

    \I__1947\ : Span4Mux_h
    port map (
            O => \N__20554\,
            I => \N__20551\
        );

    \I__1946\ : Odrv4
    port map (
            O => \N__20551\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__20548\,
            I => \N__20545\
        );

    \I__1944\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20542\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__20542\,
            I => \N__20539\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__20539\,
            I => \N__20536\
        );

    \I__1941\ : Span4Mux_v
    port map (
            O => \N__20536\,
            I => \N__20533\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__20533\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1939\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20527\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__20527\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__1937\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20521\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__20521\,
            I => \N__20518\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__20518\,
            I => \N__20515\
        );

    \I__1934\ : Odrv4
    port map (
            O => \N__20515\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__20512\,
            I => \N__20509\
        );

    \I__1932\ : InMux
    port map (
            O => \N__20509\,
            I => \N__20506\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__20506\,
            I => \N__20503\
        );

    \I__1930\ : Span4Mux_h
    port map (
            O => \N__20503\,
            I => \N__20500\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__20500\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__20497\,
            I => \N__20494\
        );

    \I__1927\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20491\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__20491\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__1925\ : InMux
    port map (
            O => \N__20488\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1924\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20482\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__20482\,
            I => \N__20479\
        );

    \I__1922\ : Span4Mux_v
    port map (
            O => \N__20479\,
            I => \N__20476\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__20476\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__20473\,
            I => \N__20470\
        );

    \I__1919\ : InMux
    port map (
            O => \N__20470\,
            I => \N__20467\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__20467\,
            I => \N__20464\
        );

    \I__1917\ : Span4Mux_h
    port map (
            O => \N__20464\,
            I => \N__20461\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__20461\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1915\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20455\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__20455\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__1913\ : InMux
    port map (
            O => \N__20452\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1912\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20446\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__20446\,
            I => \N__20443\
        );

    \I__1910\ : Span4Mux_s3_h
    port map (
            O => \N__20443\,
            I => \N__20440\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__20440\,
            I => \N__20437\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__20437\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__20434\,
            I => \N__20431\
        );

    \I__1906\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20428\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__20428\,
            I => \N__20425\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__20425\,
            I => \N__20422\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__20422\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1902\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20416\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__20416\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__1900\ : InMux
    port map (
            O => \N__20413\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1899\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20407\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__20407\,
            I => \N__20404\
        );

    \I__1897\ : Span4Mux_v
    port map (
            O => \N__20404\,
            I => \N__20401\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__20401\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__20398\,
            I => \N__20395\
        );

    \I__1894\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20392\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__20392\,
            I => \N__20389\
        );

    \I__1892\ : Span4Mux_v
    port map (
            O => \N__20389\,
            I => \N__20386\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__20386\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1890\ : InMux
    port map (
            O => \N__20383\,
            I => \N__20380\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__20380\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__1888\ : InMux
    port map (
            O => \N__20377\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1887\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20370\
        );

    \I__1886\ : InMux
    port map (
            O => \N__20373\,
            I => \N__20367\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__20370\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__20367\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1883\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20359\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__20359\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__20356\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_\
        );

    \I__1880\ : InMux
    port map (
            O => \N__20353\,
            I => \N__20349\
        );

    \I__1879\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20346\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__20349\,
            I => \N__20341\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__20346\,
            I => \N__20341\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__20341\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1875\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20333\
        );

    \I__1874\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20330\
        );

    \I__1873\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20327\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__20333\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__20330\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__20327\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__20320\,
            I => \N__20317\
        );

    \I__1868\ : InMux
    port map (
            O => \N__20317\,
            I => \N__20314\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__20314\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__1866\ : InMux
    port map (
            O => \N__20311\,
            I => \N__20308\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__20308\,
            I => \N__20304\
        );

    \I__1864\ : InMux
    port map (
            O => \N__20307\,
            I => \N__20301\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__20304\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__20301\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1861\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20293\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__20293\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__1859\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20285\
        );

    \I__1858\ : InMux
    port map (
            O => \N__20289\,
            I => \N__20280\
        );

    \I__1857\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20280\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__20285\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__20280\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__20275\,
            I => \N__20272\
        );

    \I__1853\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20268\
        );

    \I__1852\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20265\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__20268\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__20265\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1849\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20256\
        );

    \I__1848\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20253\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__20256\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__20253\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__1845\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20242\
        );

    \I__1844\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20242\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__20242\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1842\ : InMux
    port map (
            O => \N__20239\,
            I => \N__20236\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__20236\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__20233\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\
        );

    \I__1839\ : InMux
    port map (
            O => \N__20230\,
            I => \N__20226\
        );

    \I__1838\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20223\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__20226\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__20223\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__1835\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20212\
        );

    \I__1834\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20212\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__20212\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__1832\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20206\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__20206\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__20203\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\
        );

    \I__1829\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20197\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__20197\,
            I => \current_shift_inst.PI_CTRL.N_164\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__20194\,
            I => \current_shift_inst.PI_CTRL.N_164_cascade_\
        );

    \I__1826\ : InMux
    port map (
            O => \N__20191\,
            I => \N__20182\
        );

    \I__1825\ : InMux
    port map (
            O => \N__20190\,
            I => \N__20182\
        );

    \I__1824\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20182\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__20182\,
            I => \current_shift_inst.PI_CTRL.N_120\
        );

    \I__1822\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20176\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__20176\,
            I => \current_shift_inst.PI_CTRL.N_167\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__20173\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__20170\,
            I => \N__20167\
        );

    \I__1818\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20164\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__20164\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1816\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20158\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__20158\,
            I => \current_shift_inst.PI_CTRL.N_168\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__20155\,
            I => \current_shift_inst.PI_CTRL.N_27_cascade_\
        );

    \I__1813\ : InMux
    port map (
            O => \N__20152\,
            I => \N__20148\
        );

    \I__1812\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20145\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__20148\,
            I => \current_shift_inst.PI_CTRL.N_166\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__20145\,
            I => \current_shift_inst.PI_CTRL.N_166\
        );

    \I__1809\ : InMux
    port map (
            O => \N__20140\,
            I => \N__20135\
        );

    \I__1808\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20132\
        );

    \I__1807\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20129\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__20135\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__20132\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__20129\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__20122\,
            I => \N__20119\
        );

    \I__1802\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20116\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__20116\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__1800\ : InMux
    port map (
            O => \N__20113\,
            I => \N__20110\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__20110\,
            I => \N__20107\
        );

    \I__1798\ : Span4Mux_h
    port map (
            O => \N__20107\,
            I => \N__20103\
        );

    \I__1797\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20100\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__20103\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__20100\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__20095\,
            I => \N__20092\
        );

    \I__1793\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20089\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__20089\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__1791\ : InMux
    port map (
            O => \N__20086\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__1790\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20080\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__20080\,
            I => \N__20076\
        );

    \I__1788\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20073\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__20076\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__20073\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__20068\,
            I => \N__20065\
        );

    \I__1784\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20062\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__20062\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \I__1782\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20056\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__20056\,
            I => \N_34_i_i\
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__20053\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\
        );

    \I__1779\ : InMux
    port map (
            O => \N__20050\,
            I => \N__20046\
        );

    \I__1778\ : InMux
    port map (
            O => \N__20049\,
            I => \N__20043\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__20046\,
            I => \N__20040\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__20043\,
            I => pwm_duty_input_0
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__20040\,
            I => pwm_duty_input_0
        );

    \I__1774\ : InMux
    port map (
            O => \N__20035\,
            I => \N__20031\
        );

    \I__1773\ : InMux
    port map (
            O => \N__20034\,
            I => \N__20028\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__20031\,
            I => \N__20025\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__20028\,
            I => pwm_duty_input_1
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__20025\,
            I => pwm_duty_input_1
        );

    \I__1769\ : InMux
    port map (
            O => \N__20020\,
            I => \N__20016\
        );

    \I__1768\ : InMux
    port map (
            O => \N__20019\,
            I => \N__20013\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__20016\,
            I => \N__20010\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__20013\,
            I => pwm_duty_input_2
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__20010\,
            I => pwm_duty_input_2
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__20005\,
            I => \N__20002\
        );

    \I__1763\ : InMux
    port map (
            O => \N__20002\,
            I => \N__19995\
        );

    \I__1762\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19995\
        );

    \I__1761\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19992\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__19995\,
            I => pwm_duty_input_7
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__19992\,
            I => pwm_duty_input_7
        );

    \I__1758\ : InMux
    port map (
            O => \N__19987\,
            I => \N__19984\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__19984\,
            I => \N__19979\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19974\
        );

    \I__1755\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19974\
        );

    \I__1754\ : Span4Mux_v
    port map (
            O => \N__19979\,
            I => \N__19971\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__19974\,
            I => pwm_duty_input_5
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__19971\,
            I => pwm_duty_input_5
        );

    \I__1751\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19961\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19965\,
            I => \N__19958\
        );

    \I__1749\ : InMux
    port map (
            O => \N__19964\,
            I => \N__19955\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__19961\,
            I => \N__19952\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__19958\,
            I => pwm_duty_input_8
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__19955\,
            I => pwm_duty_input_8
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__19952\,
            I => pwm_duty_input_8
        );

    \I__1744\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19938\
        );

    \I__1743\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19938\
        );

    \I__1742\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19935\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__19938\,
            I => pwm_duty_input_9
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__19935\,
            I => pwm_duty_input_9
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__19930\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__1738\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19920\
        );

    \I__1737\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19920\
        );

    \I__1736\ : InMux
    port map (
            O => \N__19925\,
            I => \N__19917\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__19920\,
            I => pwm_duty_input_6
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__19917\,
            I => pwm_duty_input_6
        );

    \I__1733\ : InMux
    port map (
            O => \N__19912\,
            I => \N__19909\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__19909\,
            I => \N__19906\
        );

    \I__1731\ : Span4Mux_v
    port map (
            O => \N__19906\,
            I => \N__19903\
        );

    \I__1730\ : Odrv4
    port map (
            O => \N__19903\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1729\ : InMux
    port map (
            O => \N__19900\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__1728\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19894\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__19894\,
            I => \N__19891\
        );

    \I__1726\ : Span4Mux_v
    port map (
            O => \N__19891\,
            I => \N__19888\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__19888\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1724\ : InMux
    port map (
            O => \N__19885\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__1723\ : InMux
    port map (
            O => \N__19882\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__1722\ : InMux
    port map (
            O => \N__19879\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__1721\ : InMux
    port map (
            O => \N__19876\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__1720\ : InMux
    port map (
            O => \N__19873\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__1719\ : InMux
    port map (
            O => \N__19870\,
            I => \bfn_1_11_0_\
        );

    \I__1718\ : InMux
    port map (
            O => \N__19867\,
            I => \bfn_1_9_0_\
        );

    \I__1717\ : InMux
    port map (
            O => \N__19864\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__1716\ : InMux
    port map (
            O => \N__19861\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__1715\ : InMux
    port map (
            O => \N__19858\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__1714\ : InMux
    port map (
            O => \N__19855\,
            I => \N__19851\
        );

    \I__1713\ : InMux
    port map (
            O => \N__19854\,
            I => \N__19848\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__19851\,
            I => \N__19843\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__19848\,
            I => \N__19843\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__19843\,
            I => \N__19840\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__19840\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1708\ : InMux
    port map (
            O => \N__19837\,
            I => \N__19834\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__19834\,
            I => \N__19831\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__19831\,
            I => \N__19828\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__19828\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1704\ : InMux
    port map (
            O => \N__19825\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__1703\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19819\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__19819\,
            I => \N__19816\
        );

    \I__1701\ : Span4Mux_h
    port map (
            O => \N__19816\,
            I => \N__19813\
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__19813\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1699\ : InMux
    port map (
            O => \N__19810\,
            I => \N__19807\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__19807\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__1697\ : InMux
    port map (
            O => \N__19804\,
            I => \N__19801\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__19801\,
            I => \N__19798\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__19798\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1694\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19792\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__19792\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__1692\ : InMux
    port map (
            O => \N__19789\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__1691\ : InMux
    port map (
            O => \N__19786\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__1690\ : InMux
    port map (
            O => \N__19783\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__1689\ : InMux
    port map (
            O => \N__19780\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__1688\ : InMux
    port map (
            O => \N__19777\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__1687\ : InMux
    port map (
            O => \N__19774\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__1686\ : InMux
    port map (
            O => \N__19771\,
            I => \N__19768\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__19768\,
            I => \N__19765\
        );

    \I__1684\ : Span4Mux_h
    port map (
            O => \N__19765\,
            I => \N__19762\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__19762\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1682\ : InMux
    port map (
            O => \N__19759\,
            I => \N__19756\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__19756\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__1680\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19750\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__19750\,
            I => \N__19747\
        );

    \I__1678\ : Span4Mux_v
    port map (
            O => \N__19747\,
            I => \N__19744\
        );

    \I__1677\ : Odrv4
    port map (
            O => \N__19744\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1676\ : InMux
    port map (
            O => \N__19741\,
            I => \N__19738\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__19738\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__1674\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19732\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__19732\,
            I => \N__19729\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__19729\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1671\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19723\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__19723\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__1669\ : InMux
    port map (
            O => \N__19720\,
            I => \N__19717\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19714\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__19714\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1666\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19708\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__19708\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19702\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__19702\,
            I => \N__19699\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__19699\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1661\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19693\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__19693\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__1659\ : InMux
    port map (
            O => \N__19690\,
            I => \N__19687\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__19687\,
            I => \N__19684\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__19684\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1656\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19678\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__19678\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__1654\ : InMux
    port map (
            O => \N__19675\,
            I => \N__19672\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__19672\,
            I => \N__19669\
        );

    \I__1652\ : Span4Mux_h
    port map (
            O => \N__19669\,
            I => \N__19666\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__19666\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1650\ : InMux
    port map (
            O => \N__19663\,
            I => \N__19660\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__19660\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__1648\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19654\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__19654\,
            I => \N__19651\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__19651\,
            I => \N__19648\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__19648\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1644\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19642\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__19642\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_10_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_10_25_0_\
        );

    \IN_MUX_bfv_10_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_10_26_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_3_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_8_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_14_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_14_27_0_\
        );

    \IN_MUX_bfv_14_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_14_28_0_\
        );

    \IN_MUX_bfv_14_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_14_29_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_18_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_18_21_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_18_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_22_0_\
        );

    \IN_MUX_bfv_18_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_18_23_0_\
        );

    \IN_MUX_bfv_18_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_18_24_0_\
        );

    \IN_MUX_bfv_18_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_18_25_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_7\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_15\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_23\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            carryinitout => \bfn_13_13_0_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__22372\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_302_i_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__33295\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_180_i_g\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__39223\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_304_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__38086\,
            CLKHFEN => \N__38087\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__38162\,
            RGB2PWM => \N__20059\,
            RGB1 => rgb_g_wire,
            CURREN => \N__38163\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__20959\,
            RGB0PWM => \N__49790\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__24082\,
            in1 => \N__22820\,
            in2 => \N__24624\,
            in3 => \N__22743\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50278\,
            ce => 'H',
            sr => \N__49667\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__23989\,
            in1 => \N__22821\,
            in2 => \N__24625\,
            in3 => \N__22744\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50278\,
            ce => 'H',
            sr => \N__49667\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23788\,
            in2 => \_gnd_net_\,
            in3 => \N__20190\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => 'H',
            sr => \N__49674\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__24130\,
            in1 => \N__20950\,
            in2 => \N__20170\,
            in3 => \N__22742\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => 'H',
            sr => \N__49674\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__23755\,
            in1 => \N__20200\,
            in2 => \_gnd_net_\,
            in3 => \N__20152\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => 'H',
            sr => \N__49674\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20191\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23773\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => 'H',
            sr => \N__49674\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23803\,
            in2 => \_gnd_net_\,
            in3 => \N__20189\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => 'H',
            sr => \N__49674\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24601\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50276\,
            ce => 'H',
            sr => \N__49681\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__24049\,
            in1 => \N__22815\,
            in2 => \N__24616\,
            in3 => \N__22745\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50276\,
            ce => 'H',
            sr => \N__49681\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__22747\,
            in1 => \N__24608\,
            in2 => \N__22822\,
            in3 => \N__23956\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50276\,
            ce => 'H',
            sr => \N__49681\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__24019\,
            in1 => \N__22816\,
            in2 => \N__24617\,
            in3 => \N__22746\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50276\,
            ce => 'H',
            sr => \N__49681\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19759\,
            in2 => \_gnd_net_\,
            in3 => \N__19771\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19741\,
            in2 => \_gnd_net_\,
            in3 => \N__19753\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19726\,
            in2 => \_gnd_net_\,
            in3 => \N__19735\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19711\,
            in2 => \_gnd_net_\,
            in3 => \N__19720\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19705\,
            in1 => \N__19696\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19681\,
            in2 => \_gnd_net_\,
            in3 => \N__19690\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19663\,
            in2 => \_gnd_net_\,
            in3 => \N__19675\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19645\,
            in2 => \_gnd_net_\,
            in3 => \N__19657\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19810\,
            in2 => \_gnd_net_\,
            in3 => \N__19822\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19795\,
            in2 => \_gnd_net_\,
            in3 => \N__19804\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20631\,
            in2 => \_gnd_net_\,
            in3 => \N__19789\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__21290\,
            in1 => \N__19855\,
            in2 => \_gnd_net_\,
            in3 => \N__19786\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20138\,
            in2 => \_gnd_net_\,
            in3 => \N__19783\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20576\,
            in2 => \_gnd_net_\,
            in3 => \N__19780\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20373\,
            in2 => \_gnd_net_\,
            in3 => \N__19777\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20336\,
            in2 => \_gnd_net_\,
            in3 => \N__19774\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20288\,
            in2 => \_gnd_net_\,
            in3 => \N__19867\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20259\,
            in2 => \_gnd_net_\,
            in3 => \N__19864\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20229\,
            in2 => \_gnd_net_\,
            in3 => \N__19861\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19858\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20289\,
            in2 => \_gnd_net_\,
            in3 => \N__20271\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20106\,
            in2 => \_gnd_net_\,
            in3 => \N__20140\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20338\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20307\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19854\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19837\,
            in2 => \_gnd_net_\,
            in3 => \N__19825\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19912\,
            in2 => \_gnd_net_\,
            in3 => \N__19900\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19897\,
            in2 => \_gnd_net_\,
            in3 => \N__19885\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20530\,
            in2 => \_gnd_net_\,
            in3 => \N__19882\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38339\,
            in2 => \N__20497\,
            in3 => \N__19879\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20458\,
            in2 => \N__38386\,
            in3 => \N__19876\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20419\,
            in2 => \N__38387\,
            in3 => \N__19873\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20383\,
            in2 => \_gnd_net_\,
            in3 => \N__19870\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20848\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20812\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20776\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20737\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20701\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20677\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20656\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21097\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21076\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21052\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20986\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20086\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20079\,
            in1 => \N__21033\,
            in2 => \_gnd_net_\,
            in3 => \N__21601\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__20083\,
            in1 => \N__21037\,
            in2 => \N__20068\,
            in3 => \N__21568\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_0_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22333\,
            in2 => \_gnd_net_\,
            in3 => \N__49789\,
            lcout => \N_34_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19983\,
            in1 => \N__19927\,
            in2 => \N__20005\,
            in3 => \N__19945\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__19965\,
            in1 => \N__20935\,
            in2 => \N__20053\,
            in3 => \N__20901\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20049\,
            in1 => \N__20034\,
            in2 => \_gnd_net_\,
            in3 => \N__20019\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20001\,
            in2 => \_gnd_net_\,
            in3 => \N__19982\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__19964\,
            in1 => \N__19944\,
            in2 => \N__19930\,
            in3 => \N__19926\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__24136\,
            in1 => \N__21181\,
            in2 => \N__24614\,
            in3 => \N__22813\,
            lcout => \current_shift_inst.PI_CTRL.N_164\,
            ltout => \current_shift_inst.PI_CTRL.N_164_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__23751\,
            in1 => \N__20179\,
            in2 => \N__20194\,
            in3 => \N__20151\,
            lcout => \current_shift_inst.PI_CTRL.N_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__24593\,
            in1 => \N__21180\,
            in2 => \_gnd_net_\,
            in3 => \N__22812\,
            lcout => \current_shift_inst.PI_CTRL.N_167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24131\,
            in2 => \_gnd_net_\,
            in3 => \N__23744\,
            lcout => \current_shift_inst.PI_CTRL.N_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24077\,
            in2 => \_gnd_net_\,
            in3 => \N__23985\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23955\,
            in1 => \N__24018\,
            in2 => \N__20173\,
            in3 => \N__24048\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => \current_shift_inst.PI_CTRL.N_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__24600\,
            in1 => \N__20161\,
            in2 => \N__20155\,
            in3 => \N__22726\,
            lcout => \current_shift_inst.PI_CTRL.N_166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__21295\,
            in1 => \N__20139\,
            in2 => \N__20122\,
            in3 => \N__20113\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__20581\,
            in1 => \N__20596\,
            in2 => \N__20095\,
            in3 => \N__21297\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20374\,
            in2 => \_gnd_net_\,
            in3 => \N__20352\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__21296\,
            in1 => \N__20362\,
            in2 => \N__20356\,
            in3 => \N__20353\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__21298\,
            in1 => \N__20337\,
            in2 => \N__20320\,
            in3 => \N__20311\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__20296\,
            in1 => \N__20290\,
            in2 => \N__20275\,
            in3 => \N__21292\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20247\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20248\,
            in1 => \N__20239\,
            in2 => \N__20233\,
            in3 => \N__21293\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20230\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20217\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20218\,
            in1 => \N__20209\,
            in2 => \N__20203\,
            in3 => \N__21294\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20632\,
            in2 => \_gnd_net_\,
            in3 => \N__20619\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20620\,
            in1 => \N__20605\,
            in2 => \N__20599\,
            in3 => \N__21291\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20580\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20592\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20560\,
            in2 => \N__20548\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20524\,
            in2 => \N__20512\,
            in3 => \N__20488\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20485\,
            in2 => \N__20473\,
            in3 => \N__20452\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20449\,
            in2 => \N__20434\,
            in3 => \N__20413\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20410\,
            in2 => \N__20398\,
            in3 => \N__20377\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20875\,
            in2 => \N__20863\,
            in3 => \N__20842\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20839\,
            in2 => \N__20827\,
            in3 => \N__20806\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20803\,
            in2 => \N__20791\,
            in3 => \N__20770\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20767\,
            in2 => \N__20752\,
            in3 => \N__20731\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20728\,
            in2 => \N__20716\,
            in3 => \N__20695\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21018\,
            in2 => \N__20692\,
            in3 => \N__20671\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20668\,
            in2 => \N__21034\,
            in3 => \N__20650\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21022\,
            in2 => \N__20647\,
            in3 => \N__21091\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21088\,
            in2 => \N__21035\,
            in3 => \N__21070\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21026\,
            in2 => \N__21067\,
            in3 => \N__21046\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21043\,
            in2 => \N__21036\,
            in3 => \N__20980\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20977\,
            in2 => \N__20971\,
            in3 => \N__20962\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22332\,
            in2 => \_gnd_net_\,
            in3 => \N__49788\,
            lcout => \rgb_drv_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__24135\,
            in1 => \N__21179\,
            in2 => \N__24615\,
            in3 => \N__22814\,
            lcout => \current_shift_inst.PI_CTRL.N_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_3_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111011"
        )
    port map (
            in0 => \N__20941\,
            in1 => \N__20934\,
            in2 => \N__20911\,
            in3 => \N__20900\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23984\,
            in2 => \_gnd_net_\,
            in3 => \N__24047\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__23948\,
            in1 => \N__24017\,
            in2 => \N__21184\,
            in3 => \N__24078\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21163\,
            in2 => \N__21304\,
            in3 => \N__21303\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_8_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21157\,
            in2 => \_gnd_net_\,
            in3 => \N__21148\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21145\,
            in2 => \_gnd_net_\,
            in3 => \N__21139\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21136\,
            in2 => \_gnd_net_\,
            in3 => \N__21130\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21127\,
            in2 => \_gnd_net_\,
            in3 => \N__21121\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21118\,
            in2 => \_gnd_net_\,
            in3 => \N__21112\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21109\,
            in2 => \_gnd_net_\,
            in3 => \N__21100\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21334\,
            in2 => \_gnd_net_\,
            in3 => \N__21328\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21325\,
            in3 => \N__21316\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__21313\,
            in1 => \N__21302\,
            in2 => \N__21235\,
            in3 => \N__21220\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__21624\,
            in1 => \N__21413\,
            in2 => \N__21217\,
            in3 => \N__21462\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50264\,
            ce => 'H',
            sr => \N__49693\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__21461\,
            in1 => \N__21208\,
            in2 => \N__21418\,
            in3 => \N__21625\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50264\,
            ce => 'H',
            sr => \N__49693\
        );

    \pwm_generator_inst.threshold_8_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21202\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50260\,
            ce => 'H',
            sr => \N__49701\
        );

    \CONSTANT_ONE_LUT4_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__21620\,
            in1 => \N__21395\,
            in2 => \N__21463\,
            in3 => \N__21196\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \N__49675\
        );

    \pwm_generator_inst.threshold_4_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21190\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \N__49675\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__21394\,
            in1 => \N__21444\,
            in2 => \N__21628\,
            in3 => \N__21664\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \N__49675\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__21610\,
            in1 => \N__21464\,
            in2 => \N__21414\,
            in3 => \N__21658\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50265\,
            ce => 'H',
            sr => \N__49682\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100011011"
        )
    port map (
            in0 => \N__21613\,
            in1 => \N__21469\,
            in2 => \N__21417\,
            in3 => \N__21652\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50265\,
            ce => 'H',
            sr => \N__49682\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110101"
        )
    port map (
            in0 => \N__21468\,
            in1 => \N__21406\,
            in2 => \N__21627\,
            in3 => \N__21646\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50265\,
            ce => 'H',
            sr => \N__49682\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100011011"
        )
    port map (
            in0 => \N__21611\,
            in1 => \N__21465\,
            in2 => \N__21415\,
            in3 => \N__21640\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50265\,
            ce => 'H',
            sr => \N__49682\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__21467\,
            in1 => \N__21405\,
            in2 => \N__21626\,
            in3 => \N__21634\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50265\,
            ce => 'H',
            sr => \N__49682\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__21612\,
            in1 => \N__21466\,
            in2 => \N__21416\,
            in3 => \N__21352\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50265\,
            ce => 'H',
            sr => \N__49682\
        );

    \pwm_generator_inst.threshold_1_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21346\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50261\,
            ce => 'H',
            sr => \N__49688\
        );

    \pwm_generator_inst.threshold_6_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21340\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50261\,
            ce => 'H',
            sr => \N__49688\
        );

    \pwm_generator_inst.threshold_7_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21712\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50261\,
            ce => 'H',
            sr => \N__49688\
        );

    \pwm_generator_inst.threshold_5_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21706\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50254\,
            ce => 'H',
            sr => \N__49694\
        );

    \pwm_generator_inst.threshold_2_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21697\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50254\,
            ce => 'H',
            sr => \N__49694\
        );

    \pwm_generator_inst.threshold_3_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21688\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50254\,
            ce => 'H',
            sr => \N__49694\
        );

    \pwm_generator_inst.threshold_9_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21679\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50254\,
            ce => 'H',
            sr => \N__49694\
        );

    \phase_controller_inst1.state_1_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__22591\,
            in1 => \N__22625\,
            in2 => \N__26051\,
            in3 => \N__23884\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50215\,
            ce => 'H',
            sr => \N__49732\
        );

    \pwm_generator_inst.counter_0_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21985\,
            in1 => \N__21923\,
            in2 => \_gnd_net_\,
            in3 => \N__21673\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49668\
        );

    \pwm_generator_inst.counter_1_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21981\,
            in1 => \N__21884\,
            in2 => \_gnd_net_\,
            in3 => \N__21670\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49668\
        );

    \pwm_generator_inst.counter_2_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21986\,
            in1 => \N__21845\,
            in2 => \_gnd_net_\,
            in3 => \N__21667\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49668\
        );

    \pwm_generator_inst.counter_3_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21982\,
            in1 => \N__21809\,
            in2 => \_gnd_net_\,
            in3 => \N__21739\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49668\
        );

    \pwm_generator_inst.counter_4_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21987\,
            in1 => \N__21764\,
            in2 => \_gnd_net_\,
            in3 => \N__21736\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49668\
        );

    \pwm_generator_inst.counter_5_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21983\,
            in1 => \N__22196\,
            in2 => \_gnd_net_\,
            in3 => \N__21733\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49668\
        );

    \pwm_generator_inst.counter_6_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21988\,
            in1 => \N__22169\,
            in2 => \_gnd_net_\,
            in3 => \N__21730\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49668\
        );

    \pwm_generator_inst.counter_7_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21984\,
            in1 => \N__22124\,
            in2 => \_gnd_net_\,
            in3 => \N__21727\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__50266\,
            ce => 'H',
            sr => \N__49668\
        );

    \pwm_generator_inst.counter_8_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21980\,
            in1 => \N__22079\,
            in2 => \_gnd_net_\,
            in3 => \N__21724\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__50262\,
            ce => 'H',
            sr => \N__49676\
        );

    \pwm_generator_inst.counter_9_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__22041\,
            in1 => \N__21979\,
            in2 => \_gnd_net_\,
            in3 => \N__21721\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => 'H',
            sr => \N__49676\
        );

    \pwm_generator_inst.threshold_0_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21718\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => 'H',
            sr => \N__49676\
        );

    \pwm_generator_inst.counter_RNITBL3_9_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22198\,
            in1 => \N__22040\,
            in2 => \_gnd_net_\,
            in3 => \N__22080\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_6_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22126\,
            in1 => \N__22171\,
            in2 => \N__21991\,
            in3 => \N__21943\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIRPD2_0_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21885\,
            in2 => \_gnd_net_\,
            in3 => \N__21924\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_2_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__21847\,
            in1 => \N__21766\,
            in2 => \N__21946\,
            in3 => \N__21811\,
            lcout => \pwm_generator_inst.un1_counterlt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21901\,
            in2 => \N__21937\,
            in3 => \N__21925\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21862\,
            in2 => \N__21895\,
            in3 => \N__21886\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21826\,
            in2 => \N__21856\,
            in3 => \N__21846\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21790\,
            in2 => \N__21820\,
            in3 => \N__21810\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21745\,
            in2 => \N__21781\,
            in3 => \N__21765\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22177\,
            in2 => \N__22207\,
            in3 => \N__22197\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22170\,
            in1 => \N__22141\,
            in2 => \N__22150\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22102\,
            in2 => \N__22135\,
            in3 => \N__22125\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22057\,
            in2 => \N__22096\,
            in3 => \N__22081\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22021\,
            in2 => \N__22051\,
            in3 => \N__22042\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22015\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50242\,
            ce => 'H',
            sr => \N__49695\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32122\,
            in2 => \_gnd_net_\,
            in3 => \N__22259\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a3_1_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22316\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25109\,
            lcout => state_ns_i_a3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_4_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22317\,
            in2 => \_gnd_net_\,
            in3 => \N__25110\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50225\,
            ce => 'H',
            sr => \N__49711\
        );

    \phase_controller_inst1.state_2_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__32120\,
            in1 => \N__22261\,
            in2 => \N__22629\,
            in3 => \N__23880\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50216\,
            ce => 'H',
            sr => \N__49719\
        );

    \phase_controller_inst1.state_3_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__22260\,
            in1 => \N__32121\,
            in2 => \N__22492\,
            in3 => \N__22276\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50216\,
            ce => 'H',
            sr => \N__49719\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26041\,
            in2 => \_gnd_net_\,
            in3 => \N__22587\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__25132\,
            in1 => \N__25324\,
            in2 => \N__22285\,
            in3 => \N__22272\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50204\,
            ce => 'H',
            sr => \N__49733\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22558\,
            in2 => \_gnd_net_\,
            in3 => \N__22537\,
            lcout => \phase_controller_inst1.state_RNI7NN7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22840\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22222\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22213\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22396\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22381\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50255\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23815\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_1_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__22470\,
            in1 => \N__28033\,
            in2 => \N__22685\,
            in3 => \N__27999\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50243\,
            ce => 'H',
            sr => \N__49669\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26386\,
            in2 => \_gnd_net_\,
            in3 => \N__30498\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_302_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22675\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22469\,
            lcout => \phase_controller_inst2.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__29907\,
            in1 => \N__25133\,
            in2 => \N__22351\,
            in3 => \N__22342\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50231\,
            ce => 'H',
            sr => \N__49683\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__29701\,
            in1 => \N__29815\,
            in2 => \N__29959\,
            in3 => \N__22417\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50226\,
            ce => 'H',
            sr => \N__49689\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__22446\,
            in1 => \N__23035\,
            in2 => \N__22900\,
            in3 => \N__29860\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50217\,
            ce => 'H',
            sr => \N__49696\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22445\,
            in2 => \_gnd_net_\,
            in3 => \N__22431\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_3_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__26095\,
            in1 => \N__25730\,
            in2 => \N__22495\,
            in3 => \N__22491\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50217\,
            ce => 'H',
            sr => \N__49696\
        );

    \phase_controller_inst2.state_0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__22471\,
            in1 => \N__22432\,
            in2 => \N__22450\,
            in3 => \N__22686\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50217\,
            ce => 'H',
            sr => \N__49696\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23050\,
            in2 => \N__24535\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24505\,
            in2 => \_gnd_net_\,
            in3 => \N__22423\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23041\,
            in2 => \N__24484\,
            in3 => \N__22420\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24460\,
            in2 => \_gnd_net_\,
            in3 => \N__22408\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24850\,
            in2 => \_gnd_net_\,
            in3 => \N__22405\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24817\,
            in3 => \N__22402\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24793\,
            in3 => \N__22399\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24769\,
            in3 => \N__22522\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24744\,
            in2 => \_gnd_net_\,
            in3 => \N__22519\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24724\,
            in2 => \_gnd_net_\,
            in3 => \N__22516\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24706\,
            in2 => \_gnd_net_\,
            in3 => \N__22513\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24688\,
            in2 => \_gnd_net_\,
            in3 => \N__22510\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24985\,
            in2 => \_gnd_net_\,
            in3 => \N__22507\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24967\,
            in2 => \_gnd_net_\,
            in3 => \N__22504\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24949\,
            in2 => \_gnd_net_\,
            in3 => \N__22501\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24927\,
            in2 => \_gnd_net_\,
            in3 => \N__22498\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24907\,
            in2 => \_gnd_net_\,
            in3 => \N__22639\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17\,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24889\,
            in2 => \_gnd_net_\,
            in3 => \N__22636\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24871\,
            in2 => \_gnd_net_\,
            in3 => \N__22633\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22630\,
            in2 => \_gnd_net_\,
            in3 => \N__23873\,
            lcout => \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__25373\,
            in1 => \N__25633\,
            in2 => \_gnd_net_\,
            in3 => \N__25515\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__25516\,
            in1 => \_gnd_net_\,
            in2 => \N__25660\,
            in3 => \N__25374\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28081\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50189\,
            ce => \N__25176\,
            sr => \N__49720\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__22557\,
            in1 => \N__25783\,
            in2 => \N__22603\,
            in3 => \N__25814\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50183\,
            ce => 'H',
            sr => \N__49727\
        );

    \phase_controller_inst1.state_0_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__22580\,
            in1 => \N__22556\,
            in2 => \N__26062\,
            in3 => \N__22536\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50183\,
            ce => 'H',
            sr => \N__49727\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__25658\,
            in1 => \N__25385\,
            in2 => \N__23653\,
            in3 => \N__25551\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50183\,
            ce => 'H',
            sr => \N__49727\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__25550\,
            in1 => \N__25659\,
            in2 => \N__25427\,
            in3 => \N__22645\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50183\,
            ce => 'H',
            sr => \N__49727\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25778\,
            in1 => \N__23375\,
            in2 => \_gnd_net_\,
            in3 => \N__25808\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__25652\,
            in1 => \N__25532\,
            in2 => \N__25434\,
            in3 => \N__23503\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50178\,
            ce => 'H',
            sr => \N__49734\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__25529\,
            in1 => \N__25417\,
            in2 => \N__23479\,
            in3 => \N__25655\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50178\,
            ce => 'H',
            sr => \N__49734\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__25653\,
            in1 => \N__25533\,
            in2 => \N__25435\,
            in3 => \N__23449\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50178\,
            ce => 'H',
            sr => \N__49734\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__25530\,
            in1 => \N__25418\,
            in2 => \N__23425\,
            in3 => \N__25656\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50178\,
            ce => 'H',
            sr => \N__49734\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__25654\,
            in1 => \N__25534\,
            in2 => \N__25436\,
            in3 => \N__23707\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50178\,
            ce => 'H',
            sr => \N__49734\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__25531\,
            in1 => \N__25419\,
            in2 => \N__23683\,
            in3 => \N__25657\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50178\,
            ce => 'H',
            sr => \N__49734\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__25509\,
            in1 => \N__25641\,
            in2 => \N__25428\,
            in3 => \N__23620\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50173\,
            ce => 'H',
            sr => \N__49737\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__25637\,
            in1 => \N__25386\,
            in2 => \N__25552\,
            in3 => \N__23596\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50173\,
            ce => 'H',
            sr => \N__49737\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__25510\,
            in1 => \N__25642\,
            in2 => \N__25429\,
            in3 => \N__23569\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50173\,
            ce => 'H',
            sr => \N__49737\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__25638\,
            in1 => \N__25387\,
            in2 => \N__25553\,
            in3 => \N__23335\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50173\,
            ce => 'H',
            sr => \N__49737\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__25511\,
            in1 => \N__25643\,
            in2 => \N__25430\,
            in3 => \N__23305\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50173\,
            ce => 'H',
            sr => \N__49737\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__25639\,
            in1 => \N__25388\,
            in2 => \N__25554\,
            in3 => \N__23278\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50173\,
            ce => 'H',
            sr => \N__49737\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__25512\,
            in1 => \N__25644\,
            in2 => \N__25431\,
            in3 => \N__23563\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50173\,
            ce => 'H',
            sr => \N__49737\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__25640\,
            in1 => \N__25389\,
            in2 => \N__25555\,
            in3 => \N__23536\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50173\,
            ce => 'H',
            sr => \N__49737\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__25815\,
            in1 => \N__25631\,
            in2 => \N__25432\,
            in3 => \N__25513\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50167\,
            ce => \N__36399\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111000000"
        )
    port map (
            in0 => \N__25816\,
            in1 => \N__25632\,
            in2 => \N__25433\,
            in3 => \N__25514\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50167\,
            ce => \N__36399\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22690\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50163\,
            ce => 'H',
            sr => \N__49740\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22849\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24187\,
            in1 => \N__24208\,
            in2 => \N__24169\,
            in3 => \N__24223\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24669\,
            in2 => \_gnd_net_\,
            in3 => \N__23919\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24324\,
            in1 => \N__24649\,
            in2 => \N__22834\,
            in3 => \N__24301\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22756\,
            in1 => \N__22831\,
            in2 => \N__22825\,
            in3 => \N__22888\,
            lcout => \current_shift_inst.PI_CTRL.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24262\,
            in1 => \N__24276\,
            in2 => \N__24238\,
            in3 => \N__23904\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24277\,
            in1 => \N__24670\,
            in2 => \N__23926\,
            in3 => \N__24391\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22696\,
            in1 => \N__22867\,
            in2 => \N__22750\,
            in3 => \N__22861\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23905\,
            in1 => \N__24297\,
            in2 => \N__24325\,
            in3 => \N__24645\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24222\,
            in1 => \N__24234\,
            in2 => \N__24207\,
            in3 => \N__24261\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24343\,
            in2 => \_gnd_net_\,
            in3 => \N__24361\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24379\,
            in1 => \N__24390\,
            in2 => \N__22891\,
            in3 => \N__22882\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24435\,
            in1 => \N__24147\,
            in2 => \N__24408\,
            in3 => \N__24424\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24148\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24436\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24186\,
            in1 => \N__24165\,
            in2 => \N__22876\,
            in3 => \N__22873\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24342\,
            in1 => \N__24360\,
            in2 => \N__24409\,
            in3 => \N__22855\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24375\,
            in2 => \_gnd_net_\,
            in3 => \N__24423\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26464\,
            in2 => \_gnd_net_\,
            in3 => \N__28186\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50227\,
            ce => \N__25192\,
            sr => \N__49677\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__29696\,
            in1 => \N__29910\,
            in2 => \N__22966\,
            in3 => \N__29814\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => 'H',
            sr => \N__49684\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__29809\,
            in1 => \N__29698\,
            in2 => \N__29956\,
            in3 => \N__22951\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => 'H',
            sr => \N__49684\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__29694\,
            in1 => \N__29908\,
            in2 => \N__23017\,
            in3 => \N__29812\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => 'H',
            sr => \N__49684\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__29808\,
            in1 => \N__29697\,
            in2 => \N__29955\,
            in3 => \N__22942\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => 'H',
            sr => \N__49684\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__29811\,
            in1 => \N__29700\,
            in2 => \N__29958\,
            in3 => \N__22933\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => 'H',
            sr => \N__49684\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__29695\,
            in1 => \N__29909\,
            in2 => \N__22924\,
            in3 => \N__29813\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => 'H',
            sr => \N__49684\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__29810\,
            in1 => \N__29699\,
            in2 => \N__29957\,
            in3 => \N__22909\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50218\,
            ce => 'H',
            sr => \N__49684\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__29754\,
            in1 => \N__29927\,
            in2 => \_gnd_net_\,
            in3 => \N__29659\,
            lcout => \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__29926\,
            in1 => \N__29658\,
            in2 => \_gnd_net_\,
            in3 => \N__29753\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23033\,
            in2 => \_gnd_net_\,
            in3 => \N__29835\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29657\,
            in2 => \_gnd_net_\,
            in3 => \N__29752\,
            lcout => \phase_controller_inst2.stoper_tr.time_passed11\,
            ltout => \phase_controller_inst2.stoper_tr.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23044\,
            in3 => \N__29836\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110001101100"
        )
    port map (
            in0 => \N__23034\,
            in1 => \N__24534\,
            in2 => \N__29848\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__29651\,
            in1 => \N__29981\,
            in2 => \N__23005\,
            in3 => \N__29805\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49697\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__29802\,
            in1 => \N__29654\,
            in2 => \N__29991\,
            in3 => \N__22996\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49697\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__29652\,
            in1 => \N__29982\,
            in2 => \N__22990\,
            in3 => \N__29806\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49697\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__29803\,
            in1 => \N__29655\,
            in2 => \N__29992\,
            in3 => \N__22981\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49697\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__29653\,
            in1 => \N__29983\,
            in2 => \N__22975\,
            in3 => \N__29807\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49697\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__29804\,
            in1 => \N__29656\,
            in2 => \N__29993\,
            in3 => \N__23125\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50205\,
            ce => 'H',
            sr => \N__49697\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__29797\,
            in1 => \N__29963\,
            in2 => \N__23119\,
            in3 => \N__29691\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49702\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__29690\,
            in1 => \N__29801\,
            in2 => \N__29990\,
            in3 => \N__23110\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49702\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__29798\,
            in1 => \N__29964\,
            in2 => \N__23104\,
            in3 => \N__29692\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49702\
        );

    \phase_controller_inst1.start_timer_hc_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__23095\,
            in1 => \N__25134\,
            in2 => \N__30989\,
            in3 => \N__23083\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49702\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__29799\,
            in1 => \N__29965\,
            in2 => \N__23077\,
            in3 => \N__29693\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49702\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__29689\,
            in1 => \N__29800\,
            in2 => \N__29989\,
            in3 => \N__23068\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50196\,
            ce => 'H',
            sr => \N__49702\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23062\,
            in2 => \N__25066\,
            in3 => \N__23376\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23056\,
            in2 => \N__25027\,
            in3 => \N__23353\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23194\,
            in2 => \N__25057\,
            in3 => \N__23326\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23188\,
            in2 => \N__25219\,
            in3 => \N__23296\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23182\,
            in2 => \N__25249\,
            in3 => \N__23268\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23176\,
            in2 => \N__25231\,
            in3 => \N__23553\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25033\,
            in2 => \N__23170\,
            in3 => \N__25705\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23161\,
            in2 => \N__25264\,
            in3 => \N__25680\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23155\,
            in2 => \N__25048\,
            in3 => \N__25275\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23149\,
            in2 => \N__25201\,
            in3 => \N__23518\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23131\,
            in2 => \N__23143\,
            in3 => \N__23494\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23466\,
            in1 => \N__23251\,
            in2 => \N__25240\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23245\,
            in2 => \N__25210\,
            in3 => \N__23440\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23722\,
            in1 => \N__23239\,
            in2 => \N__25015\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23698\,
            in1 => \N__23233\,
            in2 => \N__25000\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23218\,
            in2 => \N__23227\,
            in3 => \N__23664\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23212\,
            in2 => \N__23404\,
            in3 => \N__23635\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23206\,
            in2 => \N__23395\,
            in3 => \N__23611\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23200\,
            in2 => \N__23386\,
            in3 => \N__23587\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23407\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29461\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50179\,
            ce => \N__25191\,
            sr => \N__49721\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29418\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50179\,
            ce => \N__25191\,
            sr => \N__49721\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29333\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50179\,
            ce => \N__25191\,
            sr => \N__49721\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25822\,
            in2 => \N__23377\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23349\,
            in2 => \_gnd_net_\,
            in3 => \N__23329\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25750\,
            in2 => \N__23325\,
            in3 => \N__23299\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23292\,
            in2 => \_gnd_net_\,
            in3 => \N__23272\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23269\,
            in2 => \_gnd_net_\,
            in3 => \N__23557\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23554\,
            in2 => \_gnd_net_\,
            in3 => \N__23530\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25704\,
            in2 => \_gnd_net_\,
            in3 => \N__23527\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25681\,
            in3 => \N__23524\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25282\,
            in3 => \N__23521\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23517\,
            in2 => \_gnd_net_\,
            in3 => \N__23497\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23493\,
            in2 => \_gnd_net_\,
            in3 => \N__23470\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23467\,
            in3 => \N__23443\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23439\,
            in2 => \_gnd_net_\,
            in3 => \N__23410\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23721\,
            in2 => \_gnd_net_\,
            in3 => \N__23701\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23697\,
            in2 => \_gnd_net_\,
            in3 => \N__23671\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23668\,
            in2 => \_gnd_net_\,
            in3 => \N__23638\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23634\,
            in2 => \_gnd_net_\,
            in3 => \N__23614\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23610\,
            in2 => \_gnd_net_\,
            in3 => \N__23590\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23586\,
            in2 => \_gnd_net_\,
            in3 => \N__23572\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25587\,
            in2 => \_gnd_net_\,
            in3 => \N__25476\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__30972\,
            in1 => \N__30896\,
            in2 => \_gnd_net_\,
            in3 => \N__30770\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_8_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__23864\,
            in1 => \N__28831\,
            in2 => \N__23893\,
            in3 => \N__25977\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50155\,
            ce => 'H',
            sr => \N__49741\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23848\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__27364\,
            in1 => \N__26179\,
            in2 => \N__49792\,
            in3 => \N__27397\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23824\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43873\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50251\,
            ce => 'H',
            sr => \N__49640\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39436\,
            in2 => \N__26188\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__50244\,
            ce => 'H',
            sr => \N__49647\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36530\,
            in2 => \N__26146\,
            in3 => \N__23776\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__50244\,
            ce => 'H',
            sr => \N__49647\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26128\,
            in2 => \N__39403\,
            in3 => \N__23758\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__50244\,
            ce => 'H',
            sr => \N__49647\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40882\,
            in2 => \N__28996\,
            in3 => \N__23725\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__50244\,
            ce => 'H',
            sr => \N__49647\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39360\,
            in2 => \N__26161\,
            in3 => \N__24085\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__50244\,
            ce => 'H',
            sr => \N__49647\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26152\,
            in2 => \N__43477\,
            in3 => \N__24052\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__50244\,
            ce => 'H',
            sr => \N__49647\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43535\,
            in2 => \N__26137\,
            in3 => \N__24022\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__50244\,
            ce => 'H',
            sr => \N__49647\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44202\,
            in2 => \N__28954\,
            in3 => \N__23992\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__50244\,
            ce => 'H',
            sr => \N__49647\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43636\,
            in2 => \N__26269\,
            in3 => \N__23959\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__50237\,
            ce => 'H',
            sr => \N__49652\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43591\,
            in2 => \N__26236\,
            in3 => \N__23929\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__50237\,
            ce => 'H',
            sr => \N__49652\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43801\,
            in2 => \N__27583\,
            in3 => \N__23908\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__50237\,
            ce => 'H',
            sr => \N__49652\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41739\,
            in2 => \N__27673\,
            in3 => \N__23896\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__50237\,
            ce => 'H',
            sr => \N__49652\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41670\,
            in2 => \N__26257\,
            in3 => \N__24265\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__50237\,
            ce => 'H',
            sr => \N__49652\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44139\,
            in2 => \N__26245\,
            in3 => \N__24253\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__50237\,
            ce => 'H',
            sr => \N__49652\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41523\,
            in2 => \N__24250\,
            in3 => \N__24226\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__50237\,
            ce => 'H',
            sr => \N__49652\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26122\,
            in2 => \N__36927\,
            in3 => \N__24211\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__50237\,
            ce => 'H',
            sr => \N__49652\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37116\,
            in2 => \N__27514\,
            in3 => \N__24190\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__50232\,
            ce => 'H',
            sr => \N__49656\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27604\,
            in2 => \N__41800\,
            in3 => \N__24172\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__50232\,
            ce => 'H',
            sr => \N__49656\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40206\,
            in2 => \N__26116\,
            in3 => \N__24151\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__50232\,
            ce => 'H',
            sr => \N__49656\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40149\,
            in2 => \N__27619\,
            in3 => \N__24139\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__50232\,
            ce => 'H',
            sr => \N__49656\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40269\,
            in2 => \N__27595\,
            in3 => \N__24427\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__50232\,
            ce => 'H',
            sr => \N__49656\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41458\,
            in2 => \N__27730\,
            in3 => \N__24412\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__50232\,
            ce => 'H',
            sr => \N__49656\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39491\,
            in2 => \N__27526\,
            in3 => \N__24394\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__50232\,
            ce => 'H',
            sr => \N__49656\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26224\,
            in2 => \N__44461\,
            in3 => \N__24382\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__50232\,
            ce => 'H',
            sr => \N__49656\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44573\,
            in2 => \N__27742\,
            in3 => \N__24364\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__50228\,
            ce => 'H',
            sr => \N__49662\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41344\,
            in2 => \N__27658\,
            in3 => \N__24346\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__50228\,
            ce => 'H',
            sr => \N__49662\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44653\,
            in2 => \N__26216\,
            in3 => \N__24328\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__50228\,
            ce => 'H',
            sr => \N__49662\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26207\,
            in2 => \N__36832\,
            in3 => \N__24304\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__50228\,
            ce => 'H',
            sr => \N__49662\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44521\,
            in2 => \N__26217\,
            in3 => \N__24280\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__50228\,
            ce => 'H',
            sr => \N__49662\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26211\,
            in2 => \N__39996\,
            in3 => \N__24652\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__50228\,
            ce => 'H',
            sr => \N__49662\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32191\,
            in2 => \N__26218\,
            in3 => \N__24631\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__50228\,
            ce => 'H',
            sr => \N__49662\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44913\,
            in1 => \N__26215\,
            in2 => \_gnd_net_\,
            in3 => \N__24628\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50228\,
            ce => 'H',
            sr => \N__49662\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__26680\,
            in1 => \N__26759\,
            in2 => \_gnd_net_\,
            in3 => \N__27828\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50219\,
            ce => \N__33917\,
            sr => \N__49670\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24511\,
            in2 => \N__26311\,
            in3 => \N__24524\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24490\,
            in2 => \N__26302\,
            in3 => \N__24501\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24477\,
            in1 => \N__24466\,
            in2 => \N__26281\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24442\,
            in2 => \N__26344\,
            in3 => \N__24459\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24835\,
            in2 => \N__26353\,
            in3 => \N__24846\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24799\,
            in2 => \N__24829\,
            in3 => \N__24810\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24775\,
            in2 => \N__26323\,
            in3 => \N__24786\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24762\,
            in1 => \N__24751\,
            in2 => \N__26335\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24730\,
            in2 => \N__26530\,
            in3 => \N__24745\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24712\,
            in2 => \N__26476\,
            in3 => \N__24723\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24694\,
            in2 => \N__26488\,
            in3 => \N__24705\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24676\,
            in2 => \N__26509\,
            in3 => \N__24687\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24973\,
            in2 => \N__26497\,
            in3 => \N__24984\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24955\,
            in2 => \N__26410\,
            in3 => \N__24966\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24937\,
            in2 => \N__33943\,
            in3 => \N__24948\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24913\,
            in2 => \N__26293\,
            in3 => \N__24931\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24895\,
            in2 => \N__26518\,
            in3 => \N__24906\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24888\,
            in1 => \N__24877\,
            in2 => \N__25084\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24859\,
            in2 => \N__25075\,
            in3 => \N__24870\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24853\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29419\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50197\,
            ce => \N__33925\,
            sr => \N__49690\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29334\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50197\,
            ce => \N__33925\,
            sr => \N__49690\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__26717\,
            in1 => \N__26639\,
            in2 => \N__27799\,
            in3 => \N__26555\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50190\,
            ce => \N__25189\,
            sr => \N__49698\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__26638\,
            in1 => \N__26715\,
            in2 => \N__27886\,
            in3 => \N__26577\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50190\,
            ce => \N__25189\,
            sr => \N__49698\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011110101"
        )
    port map (
            in0 => \N__26446\,
            in1 => \N__34047\,
            in2 => \N__27919\,
            in3 => \N__28108\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50190\,
            ce => \N__25189\,
            sr => \N__49698\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26716\,
            in2 => \_gnd_net_\,
            in3 => \N__27568\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50190\,
            ce => \N__25189\,
            sr => \N__49698\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__26718\,
            in1 => \N__26640\,
            in2 => \N__27856\,
            in3 => \N__26556\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50190\,
            ce => \N__25189\,
            sr => \N__49698\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__34046\,
            in1 => \N__33983\,
            in2 => \_gnd_net_\,
            in3 => \N__27775\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50190\,
            ce => \N__25189\,
            sr => \N__49698\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33984\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34048\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50190\,
            ce => \N__25189\,
            sr => \N__49698\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26731\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27715\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50184\,
            ce => \N__25190\,
            sr => \N__49703\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__26729\,
            in1 => \_gnd_net_\,
            in2 => \N__26670\,
            in3 => \N__27646\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50184\,
            ce => \N__25190\,
            sr => \N__49703\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26459\,
            in2 => \_gnd_net_\,
            in3 => \N__28210\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50184\,
            ce => \N__25190\,
            sr => \N__49703\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__26730\,
            in1 => \_gnd_net_\,
            in2 => \N__26671\,
            in3 => \N__27829\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50184\,
            ce => \N__25190\,
            sr => \N__49703\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__27949\,
            in1 => \N__26648\,
            in2 => \_gnd_net_\,
            in3 => \N__26728\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50184\,
            ce => \N__25190\,
            sr => \N__49703\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26460\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28162\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50184\,
            ce => \N__25190\,
            sr => \N__49703\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26458\,
            in2 => \_gnd_net_\,
            in3 => \N__28135\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50184\,
            ce => \N__25190\,
            sr => \N__49703\
        );

    \phase_controller_inst2.start_timer_hc_RNO_1_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26096\,
            in2 => \_gnd_net_\,
            in3 => \N__25737\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__30260\,
            in1 => \N__27961\,
            in2 => \N__25138\,
            in3 => \N__25135\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50180\,
            ce => 'H',
            sr => \N__49705\
        );

    \phase_controller_inst2.state_2_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__28000\,
            in1 => \N__25738\,
            in2 => \N__26103\,
            in3 => \N__28019\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50180\,
            ce => 'H',
            sr => \N__49705\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__30186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30447\,
            lcout => \phase_controller_inst2.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__30187\,
            in1 => \N__30261\,
            in2 => \N__28651\,
            in3 => \N__30448\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50180\,
            ce => 'H',
            sr => \N__49705\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__25661\,
            in1 => \N__25548\,
            in2 => \N__25437\,
            in3 => \N__25711\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50174\,
            ce => 'H',
            sr => \N__49712\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__25547\,
            in1 => \N__25420\,
            in2 => \N__25690\,
            in3 => \N__25663\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50174\,
            ce => 'H',
            sr => \N__49712\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__25662\,
            in1 => \N__25549\,
            in2 => \N__25438\,
            in3 => \N__25291\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50174\,
            ce => 'H',
            sr => \N__49712\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30184\,
            in1 => \N__30437\,
            in2 => \N__30308\,
            in3 => \N__26866\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50174\,
            ce => 'H',
            sr => \N__49712\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29456\,
            in1 => \N__29417\,
            in2 => \N__29335\,
            in3 => \N__28080\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30183\,
            in1 => \N__30436\,
            in2 => \N__30307\,
            in3 => \N__28285\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50174\,
            ce => 'H',
            sr => \N__49712\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__30843\,
            in1 => \N__30717\,
            in2 => \N__31077\,
            in3 => \N__25983\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50168\,
            ce => \N__36410\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__25984\,
            in1 => \N__31022\,
            in2 => \N__30757\,
            in3 => \N__30844\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50168\,
            ce => \N__36410\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25774\,
            in2 => \_gnd_net_\,
            in3 => \N__25806\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__25807\,
            in1 => \_gnd_net_\,
            in2 => \N__25782\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__30549\,
            in1 => \N__31748\,
            in2 => \N__31522\,
            in3 => \N__32983\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50164\,
            ce => \N__31594\,
            sr => \N__49728\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__31751\,
            in1 => \_gnd_net_\,
            in2 => \N__31521\,
            in3 => \N__31165\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50164\,
            ce => \N__31594\,
            sr => \N__49728\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__32839\,
            in1 => \N__31750\,
            in2 => \_gnd_net_\,
            in3 => \N__31493\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50164\,
            ce => \N__31594\,
            sr => \N__49728\
        );

    \phase_controller_inst1.stoper_hc.target_time_0_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__31747\,
            in1 => \N__30551\,
            in2 => \N__31520\,
            in3 => \N__33076\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50164\,
            ce => \N__31594\,
            sr => \N__49728\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__30550\,
            in1 => \N__31749\,
            in2 => \N__32796\,
            in3 => \N__31492\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50164\,
            ce => \N__31594\,
            sr => \N__49728\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25744\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25897\,
            in2 => \N__25906\,
            in3 => \N__27128\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25882\,
            in2 => \N__25891\,
            in3 => \N__27114\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25876\,
            in2 => \N__28924\,
            in3 => \N__27084\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25861\,
            in2 => \N__25870\,
            in3 => \N__27063\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25846\,
            in2 => \N__25855\,
            in3 => \N__27042\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25840\,
            in2 => \N__28696\,
            in3 => \N__27021\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25834\,
            in2 => \N__28684\,
            in3 => \N__27000\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25828\,
            in2 => \N__28867\,
            in3 => \N__27342\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27318\,
            in1 => \N__25954\,
            in2 => \N__30655\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25948\,
            in2 => \N__28843\,
            in3 => \N__27291\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25942\,
            in2 => \N__31768\,
            in3 => \N__27268\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27244\,
            in1 => \N__25936\,
            in2 => \N__30640\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25930\,
            in2 => \N__28897\,
            in3 => \N__27220\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25924\,
            in2 => \N__28855\,
            in3 => \N__27196\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25918\,
            in2 => \N__28909\,
            in3 => \N__27172\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25912\,
            in2 => \N__28711\,
            in3 => \N__27501\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26005\,
            in2 => \N__31609\,
            in3 => \N__27480\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25999\,
            in2 => \N__28939\,
            in3 => \N__27459\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25993\,
            in2 => \N__28882\,
            in3 => \N__27439\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25987\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28829\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25975\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__25976\,
            in1 => \_gnd_net_\,
            in2 => \N__27142\,
            in3 => \N__28830\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28828\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25974\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30794\,
            in1 => \N__30908\,
            in2 => \N__31104\,
            in3 => \N__27448\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50147\,
            ce => 'H',
            sr => \N__49742\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30904\,
            in1 => \N__30798\,
            in2 => \N__31100\,
            in3 => \N__27469\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50147\,
            ce => 'H',
            sr => \N__49742\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30792\,
            in1 => \N__30906\,
            in2 => \N__31102\,
            in3 => \N__27181\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50147\,
            ce => 'H',
            sr => \N__49742\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30903\,
            in1 => \N__30797\,
            in2 => \N__31099\,
            in3 => \N__27490\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50147\,
            ce => 'H',
            sr => \N__49742\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30793\,
            in1 => \N__30907\,
            in2 => \N__31103\,
            in3 => \N__27157\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50147\,
            ce => 'H',
            sr => \N__49742\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30901\,
            in1 => \N__30795\,
            in2 => \N__31097\,
            in3 => \N__27229\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50147\,
            ce => 'H',
            sr => \N__49742\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30791\,
            in1 => \N__30905\,
            in2 => \N__31101\,
            in3 => \N__27253\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50147\,
            ce => 'H',
            sr => \N__49742\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30902\,
            in1 => \N__30796\,
            in2 => \N__31098\,
            in3 => \N__27205\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50147\,
            ce => 'H',
            sr => \N__49742\
        );

    \phase_controller_inst2.S1_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26107\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50142\,
            ce => 'H',
            sr => \N__49745\
        );

    \phase_controller_inst1.S2_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26061\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50142\,
            ce => 'H',
            sr => \N__49745\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30909\,
            in1 => \N__30799\,
            in2 => \N__31094\,
            in3 => \N__27421\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50142\,
            ce => 'H',
            sr => \N__49745\
        );

    \delay_measurement_inst.hc_state_0_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__27359\,
            in1 => \N__26177\,
            in2 => \_gnd_net_\,
            in3 => \N__27385\,
            lcout => \delay_measurement_inst.hc_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50245\,
            ce => \N__36411\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33265\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50238\,
            ce => 'H',
            sr => \N__49628\
        );

    \delay_measurement_inst.start_timer_hc_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__27393\,
            in1 => \N__27363\,
            in2 => \_gnd_net_\,
            in3 => \N__26178\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50238\,
            ce => 'H',
            sr => \N__49628\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36205\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50233\,
            ce => 'H',
            sr => \N__49636\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36241\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50233\,
            ce => 'H',
            sr => \N__49636\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33241\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50233\,
            ce => 'H',
            sr => \N__49636\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36277\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50233\,
            ce => 'H',
            sr => \N__49636\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33451\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50233\,
            ce => 'H',
            sr => \N__49636\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36862\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50229\,
            ce => 'H',
            sr => \N__49641\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41572\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50229\,
            ce => 'H',
            sr => \N__49641\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36169\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50229\,
            ce => 'H',
            sr => \N__49641\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36570\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50229\,
            ce => 'H',
            sr => \N__49641\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36321\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50229\,
            ce => 'H',
            sr => \N__49641\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37064\,
            in2 => \_gnd_net_\,
            in3 => \N__44019\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__37199\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44018\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36642\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50209\,
            ce => 'H',
            sr => \N__49653\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36739\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50209\,
            ce => 'H',
            sr => \N__49653\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__26401\,
            in1 => \N__26385\,
            in2 => \_gnd_net_\,
            in3 => \N__30497\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50209\,
            ce => 'H',
            sr => \N__49653\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45117\,
            in1 => \N__45279\,
            in2 => \N__44917\,
            in3 => \N__40012\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50209\,
            ce => 'H',
            sr => \N__49653\
        );

    \current_shift_inst.PI_CTRL.prop_term_26_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44078\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50209\,
            ce => 'H',
            sr => \N__49653\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__26400\,
            in1 => \N__26384\,
            in2 => \_gnd_net_\,
            in3 => \N__30496\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_303_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__26750\,
            in1 => \N__26674\,
            in2 => \_gnd_net_\,
            in3 => \N__27635\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => \N__33928\,
            sr => \N__49663\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__26673\,
            in1 => \N__27941\,
            in2 => \_gnd_net_\,
            in3 => \N__26749\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => \N__33928\,
            sr => \N__49663\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26754\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27706\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => \N__33928\,
            sr => \N__49663\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26760\,
            in3 => \N__27566\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => \N__33928\,
            sr => \N__49663\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__26675\,
            in1 => \N__26755\,
            in2 => \N__27792\,
            in3 => \N__26562\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => \N__33928\,
            sr => \N__49663\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__26563\,
            in1 => \N__27848\,
            in2 => \N__26761\,
            in3 => \N__26676\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50199\,
            ce => \N__33928\,
            sr => \N__49663\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28067\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50191\,
            ce => \N__33921\,
            sr => \N__49671\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__26672\,
            in1 => \N__26732\,
            in2 => \N__27881\,
            in3 => \N__26581\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50191\,
            ce => \N__33921\,
            sr => \N__49671\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111011001111"
        )
    port map (
            in0 => \N__34025\,
            in1 => \N__27908\,
            in2 => \N__26457\,
            in3 => \N__28101\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50191\,
            ce => \N__33921\,
            sr => \N__49671\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29457\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50191\,
            ce => \N__33921\,
            sr => \N__49671\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26441\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28203\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50191\,
            ce => \N__33921\,
            sr => \N__49671\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26442\,
            in2 => \_gnd_net_\,
            in3 => \N__28154\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50191\,
            ce => \N__33921\,
            sr => \N__49671\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26440\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28179\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50191\,
            ce => \N__33921\,
            sr => \N__49671\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26439\,
            in2 => \_gnd_net_\,
            in3 => \N__28127\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50191\,
            ce => \N__33921\,
            sr => \N__49671\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__33966\,
            in1 => \N__34021\,
            in2 => \_gnd_net_\,
            in3 => \N__27765\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__27766\,
            in1 => \N__34026\,
            in2 => \_gnd_net_\,
            in3 => \N__33967\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50185\,
            ce => \N__33926\,
            sr => \N__49678\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27770\,
            in1 => \N__27642\,
            in2 => \N__34043\,
            in3 => \N__27948\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28099\,
            in2 => \_gnd_net_\,
            in3 => \N__27915\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110001"
        )
    port map (
            in0 => \N__27771\,
            in1 => \N__34045\,
            in2 => \N__26764\,
            in3 => \N__33968\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__27821\,
            in1 => \N__27711\,
            in2 => \_gnd_net_\,
            in3 => \N__27562\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__28100\,
            in1 => \_gnd_net_\,
            in2 => \N__26683\,
            in3 => \N__34044\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26614\,
            in1 => \N__26602\,
            in2 => \N__26596\,
            in3 => \N__26587\,
            lcout => \phase_controller_inst1.stoper_tr.N_248\,
            ltout => \phase_controller_inst1.stoper_tr.N_248_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__27849\,
            in1 => \_gnd_net_\,
            in2 => \N__26566\,
            in3 => \N__27882\,
            lcout => \phase_controller_inst1.stoper_tr.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26929\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26542\,
            in2 => \N__28768\,
            in3 => \N__28260\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26536\,
            in2 => \N__28738\,
            in3 => \N__28236\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28461\,
            in1 => \N__26812\,
            in2 => \N__28753\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26806\,
            in2 => \N__29587\,
            in3 => \N__28440\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28416\,
            in1 => \N__26800\,
            in2 => \N__26905\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28395\,
            in1 => \N__26794\,
            in2 => \N__26956\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26788\,
            in2 => \N__26890\,
            in3 => \N__28371\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26782\,
            in2 => \N__29548\,
            in3 => \N__28350\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26776\,
            in2 => \N__29536\,
            in3 => \N__28323\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26770\,
            in2 => \N__30463\,
            in3 => \N__28296\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26860\,
            in2 => \N__30628\,
            in3 => \N__28662\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28633\,
            in1 => \N__26854\,
            in2 => \N__29512\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26848\,
            in2 => \N__26980\,
            in3 => \N__28609\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28582\,
            in1 => \N__26842\,
            in2 => \N__26917\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26836\,
            in2 => \N__29524\,
            in3 => \N__28558\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26830\,
            in2 => \N__28723\,
            in3 => \N__28530\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26824\,
            in2 => \N__29572\,
            in3 => \N__28509\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26818\,
            in2 => \N__26941\,
            in3 => \N__28485\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26875\,
            in2 => \N__28780\,
            in3 => \N__28806\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26869\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30061\,
            in2 => \_gnd_net_\,
            in3 => \N__30019\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__30020\,
            in1 => \N__30065\,
            in2 => \_gnd_net_\,
            in3 => \N__28259\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__30239\,
            in1 => \N__30148\,
            in2 => \_gnd_net_\,
            in3 => \N__30435\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30188\,
            in1 => \N__30443\,
            in2 => \N__30323\,
            in3 => \N__28618\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50161\,
            ce => 'H',
            sr => \N__49706\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__30439\,
            in1 => \N__30291\,
            in2 => \N__28594\,
            in3 => \N__30192\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50161\,
            ce => 'H',
            sr => \N__49706\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30189\,
            in1 => \N__30444\,
            in2 => \N__30324\,
            in3 => \N__28567\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50161\,
            ce => 'H',
            sr => \N__49706\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__30440\,
            in1 => \N__30292\,
            in2 => \N__28543\,
            in3 => \N__30193\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50161\,
            ce => 'H',
            sr => \N__49706\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30190\,
            in1 => \N__30445\,
            in2 => \N__30325\,
            in3 => \N__28519\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50161\,
            ce => 'H',
            sr => \N__49706\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__30441\,
            in1 => \N__30293\,
            in2 => \N__28498\,
            in3 => \N__30194\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50161\,
            ce => 'H',
            sr => \N__49706\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30191\,
            in1 => \N__30446\,
            in2 => \N__30326\,
            in3 => \N__28474\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50161\,
            ce => 'H',
            sr => \N__49706\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__30442\,
            in1 => \N__30294\,
            in2 => \N__28792\,
            in3 => \N__30195\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50161\,
            ce => 'H',
            sr => \N__49706\
        );

    \phase_controller_inst2.stoper_hc.target_timeZ0Z_6_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__31497\,
            in1 => \N__31903\,
            in2 => \_gnd_net_\,
            in3 => \N__31740\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50157\,
            ce => \N__30595\,
            sr => \N__49713\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__31744\,
            in1 => \N__31501\,
            in2 => \_gnd_net_\,
            in3 => \N__31246\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50157\,
            ce => \N__30595\,
            sr => \N__49713\
        );

    \phase_controller_inst2.stoper_hc.target_time_0_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__30552\,
            in1 => \N__31741\,
            in2 => \N__31523\,
            in3 => \N__33075\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50157\,
            ce => \N__30595\,
            sr => \N__49713\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__31743\,
            in1 => \N__31500\,
            in2 => \_gnd_net_\,
            in3 => \N__31957\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50157\,
            ce => \N__30595\,
            sr => \N__49713\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31745\,
            in1 => \N__31502\,
            in2 => \_gnd_net_\,
            in3 => \N__31164\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50157\,
            ce => \N__30595\,
            sr => \N__49713\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__31498\,
            in1 => \N__32673\,
            in2 => \_gnd_net_\,
            in3 => \N__31746\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50157\,
            ce => \N__30595\,
            sr => \N__49713\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31742\,
            in1 => \N__31499\,
            in2 => \_gnd_net_\,
            in3 => \N__31852\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50157\,
            ce => \N__30595\,
            sr => \N__49713\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30893\,
            in1 => \N__30768\,
            in2 => \N__31096\,
            in3 => \N__27307\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50152\,
            ce => 'H',
            sr => \N__49722\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30892\,
            in1 => \N__30767\,
            in2 => \N__31095\,
            in3 => \N__26968\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50152\,
            ce => 'H',
            sr => \N__49722\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100010001100"
        )
    port map (
            in0 => \N__30759\,
            in1 => \N__27103\,
            in2 => \N__30925\,
            in3 => \N__31093\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50148\,
            ce => 'H',
            sr => \N__49729\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30899\,
            in1 => \N__30765\,
            in2 => \N__31107\,
            in3 => \N__27052\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50148\,
            ce => 'H',
            sr => \N__49729\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30762\,
            in1 => \N__31080\,
            in2 => \N__30924\,
            in3 => \N__27331\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50148\,
            ce => 'H',
            sr => \N__49729\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30897\,
            in1 => \N__30763\,
            in2 => \N__31105\,
            in3 => \N__27280\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50148\,
            ce => 'H',
            sr => \N__49729\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30761\,
            in1 => \N__31079\,
            in2 => \N__30923\,
            in3 => \N__26989\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50148\,
            ce => 'H',
            sr => \N__49729\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30900\,
            in1 => \N__30766\,
            in2 => \N__31108\,
            in3 => \N__27010\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50148\,
            ce => 'H',
            sr => \N__49729\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30760\,
            in1 => \N__31078\,
            in2 => \N__30922\,
            in3 => \N__27031\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50148\,
            ce => 'H',
            sr => \N__49729\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__30898\,
            in1 => \N__30764\,
            in2 => \N__31106\,
            in3 => \N__27073\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50148\,
            ce => 'H',
            sr => \N__49729\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27148\,
            in2 => \N__27141\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27115\,
            in2 => \_gnd_net_\,
            in3 => \N__27097\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27094\,
            in2 => \N__27088\,
            in3 => \N__27067\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27064\,
            in2 => \_gnd_net_\,
            in3 => \N__27046\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27043\,
            in2 => \_gnd_net_\,
            in3 => \N__27025\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27022\,
            in2 => \_gnd_net_\,
            in3 => \N__27004\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27001\,
            in2 => \_gnd_net_\,
            in3 => \N__26983\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27343\,
            in2 => \_gnd_net_\,
            in3 => \N__27325\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27322\,
            in2 => \_gnd_net_\,
            in3 => \N__27298\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_10_25_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27295\,
            in2 => \_gnd_net_\,
            in3 => \N__27271\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27267\,
            in2 => \_gnd_net_\,
            in3 => \N__27247\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27243\,
            in2 => \_gnd_net_\,
            in3 => \N__27223\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27219\,
            in2 => \_gnd_net_\,
            in3 => \N__27199\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27195\,
            in2 => \_gnd_net_\,
            in3 => \N__27175\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27171\,
            in2 => \_gnd_net_\,
            in3 => \N__27151\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27502\,
            in2 => \_gnd_net_\,
            in3 => \N__27484\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27481\,
            in2 => \_gnd_net_\,
            in3 => \N__27463\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_10_26_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27460\,
            in2 => \_gnd_net_\,
            in3 => \N__27442\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27438\,
            in2 => \_gnd_net_\,
            in3 => \N__27424\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_ibuf_gb_io_RNI79U7_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49787\,
            lcout => red_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC2_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27403\,
            lcout => delay_hc_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC1_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27415\,
            lcout => delay_hc_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.prev_hc_sig_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27392\,
            lcout => \delay_measurement_inst.prev_hc_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50239\,
            ce => 'H',
            sr => \N__49621\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__45067\,
            in1 => \N__45211\,
            in2 => \_gnd_net_\,
            in3 => \N__39241\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50234\,
            ce => 'H',
            sr => \N__49623\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33766\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIIOJ3_19_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36950\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36951\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50221\,
            ce => 'H',
            sr => \N__49637\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44266\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49642\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37147\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49642\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36610\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49642\
        );

    \delay_measurement_inst.delay_tr_reg_7_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__29248\,
            in1 => \N__29028\,
            in2 => \N__27567\,
            in3 => \N__37432\,
            lcout => measured_delay_tr_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49642\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36451\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49642\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36772\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49642\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__27988\,
            in1 => \N__30076\,
            in2 => \N__28045\,
            in3 => \N__30040\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50210\,
            ce => 'H',
            sr => \N__49642\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40330\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50206\,
            ce => 'H',
            sr => \N__49648\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41842\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50206\,
            ce => 'H',
            sr => \N__49648\
        );

    \delay_measurement_inst.delay_tr_reg_8_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__37404\,
            in1 => \N__29029\,
            in2 => \N__27710\,
            in3 => \N__29247\,
            lcout => measured_delay_tr_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50206\,
            ce => 'H',
            sr => \N__49648\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36487\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50206\,
            ce => 'H',
            sr => \N__49648\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45116\,
            in1 => \N__45280\,
            in2 => \N__44916\,
            in3 => \N__40039\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50206\,
            ce => 'H',
            sr => \N__49648\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41392\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50206\,
            ce => 'H',
            sr => \N__49648\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_30_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29470\,
            in1 => \N__44344\,
            in2 => \N__37756\,
            in3 => \N__33688\,
            lcout => \delay_measurement_inst.N_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_5_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__37486\,
            in1 => \N__36973\,
            in2 => \N__29054\,
            in3 => \N__29215\,
            lcout => measured_delay_tr_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50200\,
            ce => \N__29288\,
            sr => \N__49654\
        );

    \delay_measurement_inst.delay_tr_reg_esr_4_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__37485\,
            in1 => \N__36994\,
            in2 => \N__29053\,
            in3 => \N__29214\,
            lcout => measured_delay_tr_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50200\,
            ce => \N__29288\,
            sr => \N__49654\
        );

    \delay_measurement_inst.delay_tr_reg_esr_9_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000010"
        )
    port map (
            in0 => \N__29496\,
            in1 => \N__37927\,
            in2 => \N__29107\,
            in3 => \N__37371\,
            lcout => measured_delay_tr_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50192\,
            ce => \N__29287\,
            sr => \N__49660\
        );

    \delay_measurement_inst.delay_tr_reg_esr_10_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__37926\,
            in1 => \N__29497\,
            in2 => \_gnd_net_\,
            in3 => \N__37327\,
            lcout => measured_delay_tr_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50192\,
            ce => \N__29287\,
            sr => \N__49660\
        );

    \delay_measurement_inst.delay_tr_reg_ess_3_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__29213\,
            in1 => \N__37483\,
            in2 => \N__37039\,
            in3 => \N__29052\,
            lcout => measured_delay_tr_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50192\,
            ce => \N__29287\,
            sr => \N__49660\
        );

    \delay_measurement_inst.delay_tr_reg_esr_2_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__37481\,
            in1 => \N__44311\,
            in2 => \N__29055\,
            in3 => \N__29210\,
            lcout => measured_delay_tr_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50192\,
            ce => \N__29287\,
            sr => \N__49660\
        );

    \delay_measurement_inst.delay_tr_reg_esr_6_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__29211\,
            in1 => \N__29051\,
            in2 => \_gnd_net_\,
            in3 => \N__37484\,
            lcout => measured_delay_tr_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50192\,
            ce => \N__29287\,
            sr => \N__49660\
        );

    \delay_measurement_inst.delay_tr_reg_ess_1_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__37482\,
            in1 => \N__50305\,
            in2 => \N__29056\,
            in3 => \N__29212\,
            lcout => measured_delay_tr_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50192\,
            ce => \N__29287\,
            sr => \N__49660\
        );

    \delay_measurement_inst.delay_tr_reg_esr_13_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__29487\,
            in1 => \N__37910\,
            in2 => \_gnd_net_\,
            in3 => \N__37258\,
            lcout => measured_delay_tr_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50186\,
            ce => \N__29289\,
            sr => \N__49664\
        );

    \delay_measurement_inst.delay_tr_reg_esr_15_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__29375\,
            in1 => \N__29166\,
            in2 => \N__37931\,
            in3 => \N__37693\,
            lcout => measured_delay_tr_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50186\,
            ce => \N__29289\,
            sr => \N__49664\
        );

    \delay_measurement_inst.delay_tr_reg_esr_14_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__29488\,
            in1 => \N__37911\,
            in2 => \_gnd_net_\,
            in3 => \N__37738\,
            lcout => measured_delay_tr_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50186\,
            ce => \N__29289\,
            sr => \N__49664\
        );

    \delay_measurement_inst.delay_tr_reg_esr_16_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__37651\,
            in1 => \N__37912\,
            in2 => \_gnd_net_\,
            in3 => \N__29374\,
            lcout => measured_delay_tr_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50186\,
            ce => \N__29289\,
            sr => \N__49664\
        );

    \delay_measurement_inst.delay_tr_reg_esr_11_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__37908\,
            in1 => \N__29489\,
            in2 => \_gnd_net_\,
            in3 => \N__37303\,
            lcout => measured_delay_tr_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50186\,
            ce => \N__29289\,
            sr => \N__49664\
        );

    \delay_measurement_inst.delay_tr_reg_esr_12_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__37909\,
            in1 => \N__29490\,
            in2 => \_gnd_net_\,
            in3 => \N__37282\,
            lcout => measured_delay_tr_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50186\,
            ce => \N__29289\,
            sr => \N__49664\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28202\,
            in1 => \N__28178\,
            in2 => \N__28158\,
            in3 => \N__28131\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34444\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__29407\,
            in1 => \N__29443\,
            in2 => \N__29329\,
            in3 => \N__28066\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__30166\,
            in1 => \N__30309\,
            in2 => \_gnd_net_\,
            in3 => \N__30438\,
            lcout => \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28029\,
            in2 => \_gnd_net_\,
            in3 => \N__27989\,
            lcout => \phase_controller_inst2.start_timer_hc_RNO_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__30315\,
            in1 => \N__30182\,
            in2 => \N__28225\,
            in3 => \N__30429\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50170\,
            ce => 'H',
            sr => \N__49685\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30422\,
            in1 => \N__30319\,
            in2 => \N__30196\,
            in3 => \N__28450\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50170\,
            ce => 'H',
            sr => \N__49685\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__30316\,
            in1 => \N__30426\,
            in2 => \N__28429\,
            in3 => \N__30179\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50170\,
            ce => 'H',
            sr => \N__49685\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30423\,
            in1 => \N__30320\,
            in2 => \N__30197\,
            in3 => \N__28405\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50170\,
            ce => 'H',
            sr => \N__49685\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__30317\,
            in1 => \N__30427\,
            in2 => \N__28384\,
            in3 => \N__30180\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50170\,
            ce => 'H',
            sr => \N__49685\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30424\,
            in1 => \N__30321\,
            in2 => \N__30198\,
            in3 => \N__28360\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50170\,
            ce => 'H',
            sr => \N__49685\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__30318\,
            in1 => \N__30428\,
            in2 => \N__28339\,
            in3 => \N__30181\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50170\,
            ce => 'H',
            sr => \N__49685\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__30425\,
            in1 => \N__30322\,
            in2 => \N__30199\,
            in3 => \N__28312\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50170\,
            ce => 'H',
            sr => \N__49685\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28273\,
            in2 => \N__28267\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28237\,
            in2 => \_gnd_net_\,
            in3 => \N__28213\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30001\,
            in2 => \N__28465\,
            in3 => \N__28444\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28441\,
            in2 => \_gnd_net_\,
            in3 => \N__28420\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28417\,
            in2 => \_gnd_net_\,
            in3 => \N__28399\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28396\,
            in2 => \_gnd_net_\,
            in3 => \N__28375\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28372\,
            in2 => \_gnd_net_\,
            in3 => \N__28354\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28351\,
            in2 => \_gnd_net_\,
            in3 => \N__28330\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28327\,
            in2 => \_gnd_net_\,
            in3 => \N__28303\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28300\,
            in2 => \_gnd_net_\,
            in3 => \N__28276\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28669\,
            in2 => \_gnd_net_\,
            in3 => \N__28636\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28632\,
            in2 => \_gnd_net_\,
            in3 => \N__28612\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28608\,
            in2 => \_gnd_net_\,
            in3 => \N__28585\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28581\,
            in2 => \_gnd_net_\,
            in3 => \N__28561\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28557\,
            in2 => \_gnd_net_\,
            in3 => \N__28534\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28531\,
            in2 => \_gnd_net_\,
            in3 => \N__28513\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28510\,
            in2 => \_gnd_net_\,
            in3 => \N__28489\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28486\,
            in2 => \_gnd_net_\,
            in3 => \N__28468\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28807\,
            in2 => \_gnd_net_\,
            in3 => \N__28795\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__38779\,
            in1 => \N__31512\,
            in2 => \_gnd_net_\,
            in3 => \N__32731\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50153\,
            ce => \N__30612\,
            sr => \N__49707\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__30543\,
            in1 => \N__32982\,
            in2 => \N__31524\,
            in3 => \N__31666\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50153\,
            ce => \N__30612\,
            sr => \N__49707\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__30544\,
            in1 => \N__31327\,
            in2 => \N__31525\,
            in3 => \N__31668\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50153\,
            ce => \N__30612\,
            sr => \N__49707\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__31667\,
            in1 => \N__31513\,
            in2 => \N__32797\,
            in3 => \N__30545\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50153\,
            ce => \N__30612\,
            sr => \N__49707\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__31511\,
            in1 => \N__33026\,
            in2 => \_gnd_net_\,
            in3 => \N__31665\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50153\,
            ce => \N__30612\,
            sr => \N__49707\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__31507\,
            in1 => \N__33027\,
            in2 => \_gnd_net_\,
            in3 => \N__31716\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50149\,
            ce => \N__31582\,
            sr => \N__49714\
        );

    \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__31506\,
            in1 => \N__31897\,
            in2 => \_gnd_net_\,
            in3 => \N__31715\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50149\,
            ce => \N__31582\,
            sr => \N__49714\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31719\,
            in1 => \N__31510\,
            in2 => \_gnd_net_\,
            in3 => \N__32674\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50149\,
            ce => \N__31582\,
            sr => \N__49714\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__31508\,
            in1 => \N__31244\,
            in2 => \_gnd_net_\,
            in3 => \N__31717\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50149\,
            ce => \N__31582\,
            sr => \N__49714\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__31718\,
            in1 => \N__31509\,
            in2 => \N__30553\,
            in3 => \N__31325\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50149\,
            ce => \N__31582\,
            sr => \N__49714\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31738\,
            in1 => \N__31395\,
            in2 => \_gnd_net_\,
            in3 => \N__32893\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50143\,
            ce => \N__31584\,
            sr => \N__49723\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__31851\,
            in1 => \_gnd_net_\,
            in2 => \N__31440\,
            in3 => \N__31736\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50143\,
            ce => \N__31584\,
            sr => \N__49723\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__38778\,
            in1 => \N__31394\,
            in2 => \_gnd_net_\,
            in3 => \N__32730\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50143\,
            ce => \N__31584\,
            sr => \N__49723\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31739\,
            in1 => \N__31396\,
            in2 => \_gnd_net_\,
            in3 => \N__32947\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50143\,
            ce => \N__31584\,
            sr => \N__49723\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011110101"
        )
    port map (
            in0 => \N__31737\,
            in1 => \_gnd_net_\,
            in2 => \N__31953\,
            in3 => \N__31400\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50143\,
            ce => \N__31584\,
            sr => \N__49723\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__31393\,
            in1 => \N__31551\,
            in2 => \_gnd_net_\,
            in3 => \N__31735\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50143\,
            ce => \N__31584\,
            sr => \N__49723\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30758\,
            in2 => \_gnd_net_\,
            in3 => \N__30894\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_26_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__31782\,
            in1 => \N__41213\,
            in2 => \_gnd_net_\,
            in3 => \N__41046\,
            lcout => measured_delay_hc_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50129\,
            ce => 'H',
            sr => \N__49743\
        );

    \phase_controller_inst1.S1_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32155\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50128\,
            ce => 'H',
            sr => \N__49746\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44201\,
            in1 => \N__43527\,
            in2 => \N__43589\,
            in3 => \N__43470\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__43632\,
            in1 => \N__39343\,
            in2 => \N__28978\,
            in3 => \N__40877\,
            lcout => \current_shift_inst.PI_CTRL.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFI5U3_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43797\,
            in1 => \N__40205\,
            in2 => \N__32059\,
            in3 => \N__28975\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44652\,
            in1 => \N__41339\,
            in2 => \N__44520\,
            in3 => \N__41446\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNINKHC1_30_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36820\,
            in1 => \N__29071\,
            in2 => \N__32212\,
            in3 => \N__29080\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29140\,
            in1 => \N__28969\,
            in2 => \N__28963\,
            in3 => \N__28960\,
            lcout => \current_shift_inst.PI_CTRL.N_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36678\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50220\,
            ce => 'H',
            sr => \N__49624\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000110101111"
        )
    port map (
            in0 => \N__45237\,
            in1 => \N__45064\,
            in2 => \N__44922\,
            in3 => \N__39562\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50220\,
            ce => 'H',
            sr => \N__49624\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45060\,
            in1 => \N__45238\,
            in2 => \N__44918\,
            in3 => \N__39784\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50220\,
            ce => 'H',
            sr => \N__49624\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011111110"
        )
    port map (
            in0 => \N__45235\,
            in1 => \N__45062\,
            in2 => \N__44920\,
            in3 => \N__39769\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50220\,
            ce => 'H',
            sr => \N__49624\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45061\,
            in1 => \N__45239\,
            in2 => \N__44919\,
            in3 => \N__39736\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50220\,
            ce => 'H',
            sr => \N__49624\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011111110"
        )
    port map (
            in0 => \N__45236\,
            in1 => \N__45063\,
            in2 => \N__44921\,
            in3 => \N__39706\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50220\,
            ce => 'H',
            sr => \N__49624\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33421\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50220\,
            ce => 'H',
            sr => \N__49624\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI758M_30_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41515\,
            in1 => \N__37099\,
            in2 => \N__32211\,
            in3 => \N__44119\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41799\,
            in1 => \N__36907\,
            in2 => \N__41740\,
            in3 => \N__40259\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIKFFC1_21_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__39478\,
            in1 => \N__41454\,
            in2 => \N__28984\,
            in3 => \N__29002\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID8UD2_28_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__44513\,
            in1 => \N__29062\,
            in2 => \N__28981\,
            in3 => \N__41663\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIC35V7_28_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32047\,
            in1 => \N__29146\,
            in2 => \N__29089\,
            in3 => \N__29086\,
            lcout => \current_shift_inst.PI_CTRL.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI203B_12_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41514\,
            in2 => \_gnd_net_\,
            in3 => \N__41662\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFD8M_29_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44454\,
            in1 => \N__37098\,
            in2 => \N__44126\,
            in3 => \N__39985\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIIIAM_24_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41340\,
            in1 => \N__44650\,
            in2 => \N__36819\,
            in3 => \N__44562\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111110"
        )
    port map (
            in0 => \N__29170\,
            in1 => \N__29116\,
            in2 => \N__37936\,
            in3 => \N__29383\,
            lcout => \delay_measurement_inst.N_267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__37369\,
            in1 => \N__37474\,
            in2 => \N__50304\,
            in3 => \N__37035\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDB3B_18_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40141\,
            in2 => \_gnd_net_\,
            in3 => \N__40195\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36911\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34135\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI99AM_29_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44443\,
            in1 => \N__43789\,
            in2 => \N__44884\,
            in3 => \N__39989\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIDKK3_23_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36725\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_19_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40142\,
            in1 => \N__44867\,
            in2 => \N__39493\,
            in3 => \N__44563\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45065\,
            in1 => \N__45222\,
            in2 => \N__44914\,
            in3 => \N__39835\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50198\,
            ce => 'H',
            sr => \N__49643\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111110010"
        )
    port map (
            in0 => \N__45066\,
            in1 => \N__40054\,
            in2 => \N__44915\,
            in3 => \N__45223\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50198\,
            ce => 'H',
            sr => \N__49643\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36972\,
            in2 => \_gnd_net_\,
            in3 => \N__36993\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_287_4\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_287_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__44303\,
            in1 => \N__29128\,
            in2 => \N__29119\,
            in3 => \N__37731\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010001"
        )
    port map (
            in0 => \N__37732\,
            in1 => \N__37695\,
            in2 => \N__37381\,
            in3 => \N__29097\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__29098\,
            in1 => \N__37380\,
            in2 => \N__37699\,
            in3 => \N__29358\,
            lcout => \delay_measurement_inst.N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37278\,
            in1 => \N__37299\,
            in2 => \N__37257\,
            in3 => \N__37323\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\,
            ltout => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__37405\,
            in1 => \N__37431\,
            in2 => \N__29260\,
            in3 => \N__29357\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__29230\,
            in1 => \N__29176\,
            in2 => \N__37935\,
            in3 => \N__29224\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__29162\,
            in1 => \N__29257\,
            in2 => \N__29251\,
            in3 => \N__29209\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i\,
            ltout => \delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_2_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29233\,
            in3 => \N__49786\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_9_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37370\,
            in1 => \N__37736\,
            in2 => \N__37694\,
            in3 => \N__37480\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_15_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37686\,
            in2 => \_gnd_net_\,
            in3 => \N__29223\,
            lcout => \delay_measurement_inst.N_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__37571\,
            in1 => \N__37031\,
            in2 => \N__37532\,
            in3 => \N__44310\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__37610\,
            in1 => \N__37646\,
            in2 => \N__29185\,
            in3 => \N__29182\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__37647\,
            in1 => \N__37533\,
            in2 => \N__37615\,
            in3 => \N__37572\,
            lcout => \delay_measurement_inst.N_265\,
            ltout => \delay_measurement_inst.N_265_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001110"
        )
    port map (
            in0 => \N__37692\,
            in1 => \N__37737\,
            in2 => \N__29500\,
            in3 => \N__29373\,
            lcout => \delay_measurement_inst.N_270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVALS_28_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__37768\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37780\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48856\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50175\,
            ce => \N__48264\,
            sr => \N__49665\
        );

    \delay_measurement_inst.delay_tr_reg_esr_17_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__37932\,
            in1 => \N__37614\,
            in2 => \_gnd_net_\,
            in3 => \N__29384\,
            lcout => measured_delay_tr_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50169\,
            ce => \N__29296\,
            sr => \N__49672\
        );

    \delay_measurement_inst.delay_tr_reg_esr_18_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__29385\,
            in1 => \N__37933\,
            in2 => \_gnd_net_\,
            in3 => \N__37573\,
            lcout => measured_delay_tr_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50169\,
            ce => \N__29296\,
            sr => \N__49672\
        );

    \delay_measurement_inst.delay_tr_reg_esr_19_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__37934\,
            in1 => \N__37534\,
            in2 => \_gnd_net_\,
            in3 => \N__29386\,
            lcout => measured_delay_tr_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50169\,
            ce => \N__29296\,
            sr => \N__49672\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__38288\,
            in1 => \N__29266\,
            in2 => \_gnd_net_\,
            in3 => \N__45364\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46528\,
            in1 => \N__47755\,
            in2 => \N__46019\,
            in3 => \N__42970\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48852\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50165\,
            ce => \N__48261\,
            sr => \N__49679\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46531\,
            in1 => \N__47517\,
            in2 => \N__46168\,
            in3 => \N__47145\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__47146\,
            in1 => \N__45921\,
            in2 => \N__47521\,
            in3 => \N__46529\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__46530\,
            in1 => \N__29557\,
            in2 => \_gnd_net_\,
            in3 => \N__47314\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45397\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46527\,
            in2 => \N__29551\,
            in3 => \N__47313\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__31479\,
            in1 => \N__32946\,
            in2 => \_gnd_net_\,
            in3 => \N__31755\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50160\,
            ce => \N__30613\,
            sr => \N__49686\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__31756\,
            in1 => \N__31482\,
            in2 => \_gnd_net_\,
            in3 => \N__32001\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50160\,
            ce => \N__30613\,
            sr => \N__49686\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31754\,
            in1 => \N__31481\,
            in2 => \_gnd_net_\,
            in3 => \N__32892\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50160\,
            ce => \N__30613\,
            sr => \N__49686\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31753\,
            in1 => \N__31480\,
            in2 => \_gnd_net_\,
            in3 => \N__31281\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50160\,
            ce => \N__30613\,
            sr => \N__49686\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__31478\,
            in1 => \N__31560\,
            in2 => \_gnd_net_\,
            in3 => \N__31752\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50160\,
            ce => \N__30613\,
            sr => \N__49686\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_0_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__30032\,
            in1 => \N__30139\,
            in2 => \N__30331\,
            in3 => \N__30390\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50156\,
            ce => \N__36409\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_1_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001001010"
        )
    port map (
            in0 => \N__30389\,
            in1 => \N__30327\,
            in2 => \N__30185\,
            in3 => \N__30033\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50156\,
            ce => \N__36409\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30075\,
            in2 => \_gnd_net_\,
            in3 => \N__30031\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_0_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__29611\,
            in1 => \N__29995\,
            in2 => \N__29733\,
            in3 => \N__29859\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50156\,
            ce => \N__36409\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_1_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000110000"
        )
    port map (
            in0 => \N__29994\,
            in1 => \N__29858\,
            in2 => \N__29734\,
            in3 => \N__29612\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50156\,
            ce => \N__36409\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__37992\,
            in1 => \N__38287\,
            in2 => \_gnd_net_\,
            in3 => \N__37845\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__31484\,
            in1 => \N__32835\,
            in2 => \_gnd_net_\,
            in3 => \N__31664\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50151\,
            ce => \N__30611\,
            sr => \N__49699\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__31663\,
            in1 => \N__31485\,
            in2 => \_gnd_net_\,
            in3 => \N__31204\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50151\,
            ce => \N__30611\,
            sr => \N__49699\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__31483\,
            in1 => \N__32037\,
            in2 => \_gnd_net_\,
            in3 => \N__31662\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50151\,
            ce => \N__30611\,
            sr => \N__49699\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32834\,
            in1 => \N__31318\,
            in2 => \N__31163\,
            in3 => \N__33068\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31240\,
            in1 => \N__31202\,
            in2 => \N__33139\,
            in3 => \N__33025\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101010"
        )
    port map (
            in0 => \N__32701\,
            in1 => \N__31120\,
            in2 => \N__30562\,
            in3 => \N__32891\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32890\,
            in1 => \N__31941\,
            in2 => \N__33028\,
            in3 => \N__31850\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31239\,
            in1 => \N__31203\,
            in2 => \N__30559\,
            in3 => \N__30682\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32717\,
            in1 => \N__30661\,
            in2 => \N__30556\,
            in3 => \N__38777\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlt31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30508\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto8_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000001100"
        )
    port map (
            in0 => \N__32742\,
            in1 => \N__30681\,
            in2 => \N__31901\,
            in3 => \N__30469\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlt9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto14_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101010"
        )
    port map (
            in0 => \N__31952\,
            in1 => \N__32000\,
            in2 => \N__31123\,
            in3 => \N__31114\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto13_1_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31278\,
            in1 => \N__31558\,
            in2 => \N__31849\,
            in3 => \N__32034\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__31026\,
            in1 => \N__30895\,
            in2 => \_gnd_net_\,
            in3 => \N__30769\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31279\,
            in1 => \N__31559\,
            in2 => \N__32002\,
            in3 => \N__32035\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32939\,
            in2 => \_gnd_net_\,
            in3 => \N__32656\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__32827\,
            in1 => \_gnd_net_\,
            in2 => \N__31902\,
            in3 => \N__31156\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_12_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__30670\,
            in1 => \N__31326\,
            in2 => \N__30664\,
            in3 => \N__32743\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__31391\,
            in1 => \N__31992\,
            in2 => \_gnd_net_\,
            in3 => \N__31734\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50138\,
            ce => \N__31583\,
            sr => \N__49715\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__31732\,
            in1 => \N__31280\,
            in2 => \_gnd_net_\,
            in3 => \N__31392\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50138\,
            ce => \N__31583\,
            sr => \N__49715\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__31389\,
            in1 => \N__32036\,
            in2 => \_gnd_net_\,
            in3 => \N__31731\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50138\,
            ce => \N__31583\,
            sr => \N__49715\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__31390\,
            in1 => \N__31197\,
            in2 => \_gnd_net_\,
            in3 => \N__31733\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50138\,
            ce => \N__31583\,
            sr => \N__49715\
        );

    \delay_measurement_inst.delay_hc_reg_10_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__41199\,
            in1 => \N__35578\,
            in2 => \N__31561\,
            in3 => \N__41047\,
            lcout => measured_delay_hc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50135\,
            ce => 'H',
            sr => \N__49724\
        );

    \delay_measurement_inst.delay_hc_reg_31_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__41048\,
            in1 => \N__31401\,
            in2 => \_gnd_net_\,
            in3 => \N__41203\,
            lcout => measured_delay_hc_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50135\,
            ce => 'H',
            sr => \N__49724\
        );

    \delay_measurement_inst.delay_hc_reg_3_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__35209\,
            in1 => \N__31317\,
            in2 => \N__41219\,
            in3 => \N__41049\,
            lcout => measured_delay_hc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50135\,
            ce => 'H',
            sr => \N__49724\
        );

    \delay_measurement_inst.delay_hc_reg_12_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__41017\,
            in1 => \N__35467\,
            in2 => \N__31282\,
            in3 => \N__41156\,
            lcout => measured_delay_hc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50133\,
            ce => 'H',
            sr => \N__49730\
        );

    \delay_measurement_inst.delay_hc_reg_18_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__41154\,
            in1 => \N__39052\,
            in2 => \N__31245\,
            in3 => \N__41019\,
            lcout => measured_delay_hc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50133\,
            ce => 'H',
            sr => \N__49730\
        );

    \delay_measurement_inst.delay_hc_reg_17_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011111010"
        )
    port map (
            in0 => \N__41018\,
            in1 => \N__39022\,
            in2 => \N__31201\,
            in3 => \N__41157\,
            lcout => measured_delay_hc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50133\,
            ce => 'H',
            sr => \N__49730\
        );

    \delay_measurement_inst.delay_hc_reg_5_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41020\,
            in1 => \N__31152\,
            in2 => \N__41220\,
            in3 => \N__35143\,
            lcout => measured_delay_hc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50133\,
            ce => 'H',
            sr => \N__49730\
        );

    \delay_measurement_inst.delay_hc_reg_11_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__41153\,
            in1 => \N__35521\,
            in2 => \N__32038\,
            in3 => \N__41016\,
            lcout => measured_delay_hc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50133\,
            ce => 'H',
            sr => \N__49730\
        );

    \delay_measurement_inst.delay_hc_reg_9_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__41155\,
            in1 => \N__34924\,
            in2 => \N__31996\,
            in3 => \N__41021\,
            lcout => measured_delay_hc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50133\,
            ce => 'H',
            sr => \N__49730\
        );

    \delay_measurement_inst.delay_hc_reg_24_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__40980\,
            in1 => \_gnd_net_\,
            in2 => \N__41207\,
            in3 => \N__31807\,
            lcout => measured_delay_hc_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50131\,
            ce => 'H',
            sr => \N__49735\
        );

    \delay_measurement_inst.delay_hc_reg_14_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__35356\,
            in1 => \N__41159\,
            in2 => \N__31951\,
            in3 => \N__40979\,
            lcout => measured_delay_hc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50131\,
            ce => 'H',
            sr => \N__49735\
        );

    \delay_measurement_inst.delay_hc_reg_6_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__40982\,
            in1 => \N__31879\,
            in2 => \N__41209\,
            in3 => \N__35095\,
            lcout => measured_delay_hc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50131\,
            ce => 'H',
            sr => \N__49735\
        );

    \delay_measurement_inst.delay_hc_reg_25_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__40981\,
            in1 => \_gnd_net_\,
            in2 => \N__41208\,
            in3 => \N__31795\,
            lcout => measured_delay_hc_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50131\,
            ce => 'H',
            sr => \N__49735\
        );

    \delay_measurement_inst.delay_hc_reg_13_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__35413\,
            in1 => \N__41158\,
            in2 => \N__31848\,
            in3 => \N__40978\,
            lcout => measured_delay_hc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50131\,
            ce => 'H',
            sr => \N__49735\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_1_4_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31806\,
            in1 => \N__31794\,
            in2 => \N__31783\,
            in3 => \N__32166\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35466\,
            in1 => \N__35517\,
            in2 => \N__35412\,
            in3 => \N__35577\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__33177\,
            in1 => \N__43662\,
            in2 => \_gnd_net_\,
            in3 => \N__33319\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50127\,
            ce => 'H',
            sr => \N__49739\
        );

    \delay_measurement_inst.delay_hc_reg_23_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__41212\,
            in1 => \N__32167\,
            in2 => \_gnd_net_\,
            in3 => \N__40983\,
            lcout => measured_delay_hc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50127\,
            ce => 'H',
            sr => \N__49739\
        );

    \current_shift_inst.start_timer_s1_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__32075\,
            in1 => \N__33176\,
            in2 => \_gnd_net_\,
            in3 => \N__32147\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50127\,
            ce => 'H',
            sr => \N__49739\
        );

    \current_shift_inst.stop_timer_s1_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101100001000"
        )
    port map (
            in0 => \N__33178\,
            in1 => \N__32154\,
            in2 => \N__32082\,
            in3 => \N__33318\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50126\,
            ce => 'H',
            sr => \N__49744\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33838\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50240\,
            ce => 'H',
            sr => \N__49616\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36906\,
            in1 => \N__41789\,
            in2 => \N__40270\,
            in3 => \N__41729\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__39402\,
            in1 => \N__36517\,
            in2 => \_gnd_net_\,
            in3 => \N__39432\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un1_enablelt3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010001"
        )
    port map (
            in0 => \N__39353\,
            in1 => \N__40873\,
            in2 => \N__32050\,
            in3 => \N__43495\,
            lcout => \current_shift_inst.PI_CTRL.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36677\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36233\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36269\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36197\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32201\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36560\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36161\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIFLJ3_16_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36764\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36479\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36602\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36638\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36311\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIEKJ3_15_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36854\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32248\,
            in2 => \_gnd_net_\,
            in3 => \N__33834\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33628\,
            in2 => \_gnd_net_\,
            in3 => \N__32242\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__50211\,
            ce => 'H',
            sr => \N__49629\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33862\,
            in2 => \_gnd_net_\,
            in3 => \N__32239\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__50211\,
            ce => 'H',
            sr => \N__49629\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33727\,
            in3 => \N__32236\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__50211\,
            ce => 'H',
            sr => \N__49629\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32233\,
            in2 => \_gnd_net_\,
            in3 => \N__32221\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__50211\,
            ce => 'H',
            sr => \N__49629\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33706\,
            in2 => \_gnd_net_\,
            in3 => \N__32218\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__50211\,
            ce => 'H',
            sr => \N__49629\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32356\,
            in2 => \_gnd_net_\,
            in3 => \N__32215\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__50211\,
            ce => 'H',
            sr => \N__49629\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33592\,
            in2 => \_gnd_net_\,
            in3 => \N__32281\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__50211\,
            ce => 'H',
            sr => \N__49629\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33748\,
            in2 => \_gnd_net_\,
            in3 => \N__32278\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__50207\,
            ce => 'H',
            sr => \N__49638\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32275\,
            in2 => \_gnd_net_\,
            in3 => \N__32269\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__50207\,
            ce => 'H',
            sr => \N__49638\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33742\,
            in2 => \_gnd_net_\,
            in3 => \N__32266\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__50207\,
            ce => 'H',
            sr => \N__49638\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33652\,
            in2 => \_gnd_net_\,
            in3 => \N__32263\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__50207\,
            ce => 'H',
            sr => \N__49638\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33697\,
            in2 => \_gnd_net_\,
            in3 => \N__32260\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__50207\,
            ce => 'H',
            sr => \N__49638\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33664\,
            in2 => \_gnd_net_\,
            in3 => \N__32257\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__50207\,
            ce => 'H',
            sr => \N__49638\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33715\,
            in2 => \_gnd_net_\,
            in3 => \N__32254\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            clk => \N__50207\,
            ce => 'H',
            sr => \N__49638\
        );

    \current_shift_inst.PI_CTRL.error_control_15_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34060\,
            in2 => \_gnd_net_\,
            in3 => \N__32251\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            clk => \N__50207\,
            ce => 'H',
            sr => \N__49638\
        );

    \current_shift_inst.PI_CTRL.error_control_16_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33658\,
            in2 => \_gnd_net_\,
            in3 => \N__32320\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_16\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            clk => \N__50201\,
            ce => 'H',
            sr => \N__49644\
        );

    \current_shift_inst.PI_CTRL.error_control_17_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33277\,
            in2 => \_gnd_net_\,
            in3 => \N__32317\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            clk => \N__50201\,
            ce => 'H',
            sr => \N__49644\
        );

    \current_shift_inst.PI_CTRL.error_control_18_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33736\,
            in3 => \N__32314\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            clk => \N__50201\,
            ce => 'H',
            sr => \N__49644\
        );

    \current_shift_inst.PI_CTRL.error_control_19_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33676\,
            in2 => \_gnd_net_\,
            in3 => \N__32311\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            clk => \N__50201\,
            ce => 'H',
            sr => \N__49644\
        );

    \current_shift_inst.PI_CTRL.error_control_20_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33619\,
            in2 => \_gnd_net_\,
            in3 => \N__32308\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            clk => \N__50201\,
            ce => 'H',
            sr => \N__49644\
        );

    \current_shift_inst.PI_CTRL.error_control_21_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32329\,
            in2 => \_gnd_net_\,
            in3 => \N__32305\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            clk => \N__50201\,
            ce => 'H',
            sr => \N__49644\
        );

    \current_shift_inst.PI_CTRL.error_control_22_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32302\,
            in2 => \_gnd_net_\,
            in3 => \N__32290\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            clk => \N__50201\,
            ce => 'H',
            sr => \N__49644\
        );

    \current_shift_inst.PI_CTRL.error_control_23_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33850\,
            in2 => \_gnd_net_\,
            in3 => \N__32287\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            clk => \N__50201\,
            ce => 'H',
            sr => \N__49644\
        );

    \current_shift_inst.PI_CTRL.error_control_24_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32335\,
            in2 => \_gnd_net_\,
            in3 => \N__32284\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_24\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            clk => \N__50193\,
            ce => 'H',
            sr => \N__49649\
        );

    \current_shift_inst.PI_CTRL.error_control_25_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32341\,
            in2 => \_gnd_net_\,
            in3 => \N__32347\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            clk => \N__50193\,
            ce => 'H',
            sr => \N__49649\
        );

    \current_shift_inst.PI_CTRL.error_control_26_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34387\,
            in2 => \_gnd_net_\,
            in3 => \N__32344\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50193\,
            ce => 'H',
            sr => \N__49649\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34386\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38614\,
            in1 => \N__32554\,
            in2 => \_gnd_net_\,
            in3 => \N__46993\,
            lcout => \current_shift_inst.control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46744\,
            in1 => \N__48190\,
            in2 => \N__46341\,
            in3 => \N__42819\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__32488\,
            in1 => \N__38557\,
            in2 => \_gnd_net_\,
            in3 => \N__46994\,
            lcout => \current_shift_inst.control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46743\,
            in1 => \N__47590\,
            in2 => \N__46340\,
            in3 => \N__42880\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46026\,
            in1 => \N__46745\,
            in2 => \N__48586\,
            in3 => \N__43060\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__46995\,
            in1 => \N__38503\,
            in2 => \_gnd_net_\,
            in3 => \N__32635\,
            lcout => \current_shift_inst.control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38485\,
            in1 => \N__32620\,
            in2 => \_gnd_net_\,
            in3 => \N__46973\,
            lcout => \current_shift_inst.control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__46974\,
            in1 => \N__38734\,
            in2 => \_gnd_net_\,
            in3 => \N__32608\,
            lcout => \current_shift_inst.control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__32371\,
            in1 => \N__38419\,
            in2 => \_gnd_net_\,
            in3 => \N__46969\,
            lcout => \current_shift_inst.control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__47905\,
            in1 => \N__42558\,
            in2 => \N__46228\,
            in3 => \N__46707\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38593\,
            in1 => \N__32521\,
            in2 => \_gnd_net_\,
            in3 => \N__46970\,
            lcout => \current_shift_inst.control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34180\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__32473\,
            in1 => \N__38539\,
            in2 => \_gnd_net_\,
            in3 => \N__46971\,
            lcout => \current_shift_inst.control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__46972\,
            in1 => \N__38521\,
            in2 => \_gnd_net_\,
            in3 => \N__32458\,
            lcout => \current_shift_inst.control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__47800\,
            in1 => \N__46006\,
            in2 => \N__46742\,
            in3 => \N__42999\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__32581\,
            in1 => \N__38701\,
            in2 => \_gnd_net_\,
            in3 => \N__46980\,
            lcout => \current_shift_inst.control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46651\,
            in1 => \N__47713\,
            in2 => \N__46217\,
            in3 => \N__42936\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__32500\,
            in1 => \N__38575\,
            in2 => \_gnd_net_\,
            in3 => \N__46979\,
            lcout => \current_shift_inst.control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46647\,
            in1 => \N__47833\,
            in2 => \N__46218\,
            in3 => \N__47407\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38449\,
            in1 => \N__32410\,
            in2 => \_gnd_net_\,
            in3 => \N__46975\,
            lcout => \current_shift_inst.control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38434\,
            in2 => \N__46992\,
            in3 => \N__32392\,
            lcout => \current_shift_inst.control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__46007\,
            in1 => \N__48235\,
            in2 => \N__46797\,
            in3 => \N__42846\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32362\,
            in2 => \N__37975\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40438\,
            in2 => \N__40417\,
            in3 => \N__37843\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37844\,
            in1 => \N__32446\,
            in2 => \N__45925\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40099\,
            in2 => \N__45928\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45547\,
            in2 => \N__45926\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32440\,
            in2 => \N__45929\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45532\,
            in2 => \N__45927\,
            in3 => \N__32431\,
            lcout => \current_shift_inst.un38_control_input_0_s0_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32428\,
            in2 => \N__45930\,
            in3 => \N__32422\,
            lcout => \current_shift_inst.un38_control_input_0_s0_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32419\,
            in2 => \N__45991\,
            in3 => \N__32401\,
            lcout => \current_shift_inst.un38_control_input_0_s0_8\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32398\,
            in2 => \N__45995\,
            in3 => \N__32383\,
            lcout => \current_shift_inst.un38_control_input_0_s0_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32380\,
            in2 => \N__45992\,
            in3 => \N__32560\,
            lcout => \current_shift_inst.un38_control_input_0_s0_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47095\,
            in2 => \N__45996\,
            in3 => \N__32557\,
            lcout => \current_shift_inst.un38_control_input_0_s0_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34513\,
            in2 => \N__45993\,
            in3 => \N__32545\,
            lcout => \current_shift_inst.un38_control_input_0_s0_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32542\,
            in2 => \N__45997\,
            in3 => \N__32533\,
            lcout => \current_shift_inst.un38_control_input_0_s0_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32530\,
            in2 => \N__45994\,
            in3 => \N__32512\,
            lcout => \current_shift_inst.un38_control_input_0_s0_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32509\,
            in2 => \N__45998\,
            in3 => \N__32491\,
            lcout => \current_shift_inst.un38_control_input_0_s0_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45959\,
            in2 => \N__45487\,
            in3 => \N__32476\,
            lcout => \current_shift_inst.un38_control_input_0_s0_16\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43351\,
            in2 => \N__46208\,
            in3 => \N__32461\,
            lcout => \current_shift_inst.un38_control_input_0_s0_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45963\,
            in2 => \N__34507\,
            in3 => \N__32449\,
            lcout => \current_shift_inst.un38_control_input_0_s0_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40591\,
            in2 => \N__46209\,
            in3 => \N__32623\,
            lcout => \current_shift_inst.un38_control_input_0_s0_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45967\,
            in2 => \N__40681\,
            in3 => \N__32611\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34483\,
            in2 => \N__46210\,
            in3 => \N__32599\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45971\,
            in2 => \N__32596\,
            in3 => \N__32584\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45999\,
            in2 => \N__43150\,
            in3 => \N__32572\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34600\,
            in2 => \N__46211\,
            in3 => \N__32569\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43681\,
            in2 => \N__46215\,
            in3 => \N__32566\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34606\,
            in2 => \N__46212\,
            in3 => \N__32563\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43300\,
            in2 => \N__46216\,
            in3 => \N__32758\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34612\,
            in2 => \N__46213\,
            in3 => \N__32755\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45981\,
            in2 => \N__40711\,
            in3 => \N__32752\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40783\,
            in2 => \N__46214\,
            in3 => \N__32749\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_0_25_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__45457\,
            in1 => \N__39064\,
            in2 => \N__46996\,
            in3 => \N__32746\,
            lcout => \current_shift_inst.control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto5_2_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32778\,
            in2 => \_gnd_net_\,
            in3 => \N__32974\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33042\,
            in1 => \N__32690\,
            in2 => \N__33135\,
            in3 => \N__32911\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_1_6_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__32910\,
            in1 => \N__33041\,
            in2 => \N__32692\,
            in3 => \N__38776\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_22_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__41185\,
            in1 => \N__32691\,
            in2 => \_gnd_net_\,
            in3 => \N__41038\,
            lcout => measured_delay_hc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50144\,
            ce => 'H',
            sr => \N__49708\
        );

    \delay_measurement_inst.delay_hc_reg_7_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__41039\,
            in1 => \N__41186\,
            in2 => \N__32672\,
            in3 => \N__35044\,
            lcout => measured_delay_hc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50144\,
            ce => 'H',
            sr => \N__49708\
        );

    \delay_measurement_inst.delay_hc_reg_0_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__41183\,
            in1 => \N__33067\,
            in2 => \_gnd_net_\,
            in3 => \N__41036\,
            lcout => measured_delay_hc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50144\,
            ce => 'H',
            sr => \N__49708\
        );

    \delay_measurement_inst.delay_hc_reg_20_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__41184\,
            in1 => \N__33043\,
            in2 => \_gnd_net_\,
            in3 => \N__41037\,
            lcout => measured_delay_hc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50144\,
            ce => 'H',
            sr => \N__49708\
        );

    \delay_measurement_inst.delay_hc_reg_16_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__41195\,
            in1 => \N__38992\,
            in2 => \N__33021\,
            in3 => \N__41032\,
            lcout => measured_delay_hc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50139\,
            ce => 'H',
            sr => \N__49716\
        );

    \delay_measurement_inst.delay_hc_reg_1_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__41033\,
            in1 => \N__41197\,
            in2 => \N__32981\,
            in3 => \N__38881\,
            lcout => measured_delay_hc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50139\,
            ce => 'H',
            sr => \N__49716\
        );

    \delay_measurement_inst.delay_hc_reg_8_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__41196\,
            in1 => \N__32938\,
            in2 => \N__34987\,
            in3 => \N__41035\,
            lcout => measured_delay_hc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50139\,
            ce => 'H',
            sr => \N__49716\
        );

    \delay_measurement_inst.delay_hc_reg_21_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__41034\,
            in1 => \N__32909\,
            in2 => \_gnd_net_\,
            in3 => \N__41198\,
            lcout => measured_delay_hc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50139\,
            ce => 'H',
            sr => \N__49716\
        );

    \delay_measurement_inst.delay_hc_reg_15_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__35299\,
            in1 => \N__41169\,
            in2 => \N__32889\,
            in3 => \N__41012\,
            lcout => measured_delay_hc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50136\,
            ce => 'H',
            sr => \N__49725\
        );

    \delay_measurement_inst.delay_hc_reg_4_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__41015\,
            in1 => \N__35185\,
            in2 => \N__41211\,
            in3 => \N__32823\,
            lcout => measured_delay_hc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50136\,
            ce => 'H',
            sr => \N__49725\
        );

    \delay_measurement_inst.delay_hc_reg_2_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41014\,
            in1 => \N__32777\,
            in2 => \N__41210\,
            in3 => \N__38836\,
            lcout => measured_delay_hc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50136\,
            ce => 'H',
            sr => \N__49725\
        );

    \delay_measurement_inst.delay_hc_reg_19_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__38960\,
            in1 => \N__41170\,
            in2 => \N__33134\,
            in3 => \N__41013\,
            lcout => measured_delay_hc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50136\,
            ce => 'H',
            sr => \N__49725\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64F91_1_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__35135\,
            in1 => \N__38832\,
            in2 => \_gnd_net_\,
            in3 => \N__38877\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHDUI2_3_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__35183\,
            in1 => \N__35201\,
            in2 => \N__33103\,
            in3 => \N__35089\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64AN1_6_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__35090\,
            in1 => \N__35038\,
            in2 => \N__34986\,
            in3 => \N__34912\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35402\,
            in1 => \N__38978\,
            in2 => \N__34920\,
            in3 => \N__35091\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_11_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33214\,
            in1 => \N__33094\,
            in2 => \N__33100\,
            in3 => \N__35215\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000100"
        )
    port map (
            in0 => \N__38935\,
            in1 => \N__33328\,
            in2 => \N__33097\,
            in3 => \N__33082\,
            lcout => \delay_measurement_inst.un1_elapsed_time_hc\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_17_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35136\,
            in1 => \N__39017\,
            in2 => \N__39047\,
            in3 => \N__35184\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINEU73_14_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110101"
        )
    port map (
            in0 => \N__35348\,
            in1 => \N__33088\,
            in2 => \N__33202\,
            in3 => \N__35293\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35347\,
            in1 => \N__35459\,
            in2 => \N__35298\,
            in3 => \N__35516\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI72ES3_7_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__34916\,
            in1 => \N__35039\,
            in2 => \N__34982\,
            in3 => \N__33208\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOC2D5_14_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000110011"
        )
    port map (
            in0 => \N__33198\,
            in1 => \N__35294\,
            in2 => \N__33184\,
            in3 => \N__35349\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt19_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000110011"
        )
    port map (
            in0 => \N__38934\,
            in1 => \N__35914\,
            in2 => \N__33181\,
            in3 => \N__33151\,
            lcout => \delay_measurement_inst.delay_hc_reg3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35910\,
            in1 => \N__35718\,
            in2 => \N__35797\,
            in3 => \N__35755\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__43661\,
            in1 => \N__33175\,
            in2 => \_gnd_net_\,
            in3 => \N__33317\,
            lcout => \current_shift_inst.timer_s1.N_181_i_g\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35754\,
            in2 => \_gnd_net_\,
            in3 => \N__35719\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__35796\,
            in1 => \N__33285\,
            in2 => \N__33154\,
            in3 => \N__33145\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35617\,
            in1 => \N__35647\,
            in2 => \N__36112\,
            in3 => \N__35680\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02O13_20_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33337\,
            in2 => \N__33331\,
            in3 => \N__33286\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43657\,
            in2 => \_gnd_net_\,
            in3 => \N__33316\,
            lcout => \current_shift_inst.timer_s1.N_180_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_13_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35980\,
            in1 => \N__36034\,
            in2 => \N__35929\,
            in3 => \N__36073\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41779\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34249\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39465\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43469\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33258\,
            in1 => \N__33247\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33220\,
            in2 => \_gnd_net_\,
            in3 => \N__33237\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33427\,
            in2 => \_gnd_net_\,
            in3 => \N__33450\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33403\,
            in2 => \_gnd_net_\,
            in3 => \N__33420\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33397\,
            in2 => \_gnd_net_\,
            in3 => \N__33391\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33388\,
            in3 => \N__33379\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33376\,
            in2 => \_gnd_net_\,
            in3 => \N__33370\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33367\,
            in2 => \_gnd_net_\,
            in3 => \N__33358\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33355\,
            in2 => \_gnd_net_\,
            in3 => \N__33349\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_8\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33346\,
            in2 => \_gnd_net_\,
            in3 => \N__33340\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33520\,
            in2 => \_gnd_net_\,
            in3 => \N__33514\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33511\,
            in2 => \_gnd_net_\,
            in3 => \N__33505\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33502\,
            in2 => \_gnd_net_\,
            in3 => \N__33496\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33493\,
            in2 => \_gnd_net_\,
            in3 => \N__33487\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIDHEC_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33484\,
            in2 => \_gnd_net_\,
            in3 => \N__33478\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIFKFC_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33475\,
            in2 => \_gnd_net_\,
            in3 => \N__33469\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIHNGC_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33466\,
            in2 => \_gnd_net_\,
            in3 => \N__33460\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_16\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIJQHC_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33586\,
            in2 => \_gnd_net_\,
            in3 => \N__33457\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNILTIC_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33601\,
            in2 => \_gnd_net_\,
            in3 => \N__33454\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIN0KC_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33568\,
            in2 => \_gnd_net_\,
            in3 => \N__33559\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNIGRLC_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33637\,
            in2 => \_gnd_net_\,
            in3 => \N__33556\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNI9DFD_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33646\,
            in2 => \_gnd_net_\,
            in3 => \N__33553\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIBGGD_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33577\,
            in2 => \_gnd_net_\,
            in3 => \N__33550\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIDJHD_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33547\,
            in2 => \_gnd_net_\,
            in3 => \N__33535\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIFMID_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33670\,
            in2 => \_gnd_net_\,
            in3 => \N__33532\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_24\,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIHPJD_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41365\,
            in2 => \_gnd_net_\,
            in3 => \N__33529\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37200\,
            in2 => \_gnd_net_\,
            in3 => \N__33526\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36702\,
            in2 => \_gnd_net_\,
            in3 => \N__33523\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37065\,
            in2 => \_gnd_net_\,
            in3 => \N__33613\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37172\,
            in2 => \_gnd_net_\,
            in3 => \N__33610\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37233\,
            in2 => \_gnd_net_\,
            in3 => \N__33607\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5K_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__44017\,
            in1 => \N__36831\,
            in2 => \_gnd_net_\,
            in3 => \N__33604\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIHNJ3_18_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41558\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34171\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__37232\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43981\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIGMJ3_17_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44252\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNICJK3_22_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36437\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIELK3_24_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__37174\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43980\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34315\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34267\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34090\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBIK3_21_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41828\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIAHK3_20_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37133\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33817\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34210\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34153\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34108\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34234\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33784\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34297\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34198\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34072\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9AP1_24_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37801\,
            in1 => \N__37810\,
            in2 => \N__37792\,
            in3 => \N__37819\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34222\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34279\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34042\,
            in2 => \_gnd_net_\,
            in3 => \N__33985\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50194\,
            ce => \N__33927\,
            sr => \N__49650\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33799\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34429\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_0_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34333\,
            in2 => \N__34357\,
            in3 => \N__34356\,
            lcout => \current_shift_inst.control_inputZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.control_input_1_cry_0\,
            clk => \N__50187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34540\,
            in2 => \_gnd_net_\,
            in3 => \N__33808\,
            lcout => \current_shift_inst.control_inputZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_0\,
            carryout => \current_shift_inst.control_input_1_cry_1\,
            clk => \N__50187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_2_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33805\,
            in2 => \_gnd_net_\,
            in3 => \N__33793\,
            lcout => \current_shift_inst.control_inputZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_1\,
            carryout => \current_shift_inst.control_input_1_cry_2\,
            clk => \N__50187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_3_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33790\,
            in2 => \_gnd_net_\,
            in3 => \N__33775\,
            lcout => \current_shift_inst.control_inputZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_2\,
            carryout => \current_shift_inst.control_input_1_cry_3\,
            clk => \N__50187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_4_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33772\,
            in2 => \_gnd_net_\,
            in3 => \N__33751\,
            lcout => \current_shift_inst.control_inputZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_3\,
            carryout => \current_shift_inst.control_input_1_cry_4\,
            clk => \N__50187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_5_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47020\,
            in2 => \_gnd_net_\,
            in3 => \N__34189\,
            lcout => \current_shift_inst.control_inputZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_4\,
            carryout => \current_shift_inst.control_input_1_cry_5\,
            clk => \N__50187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_6_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34186\,
            in2 => \_gnd_net_\,
            in3 => \N__34174\,
            lcout => \current_shift_inst.control_inputZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_5\,
            carryout => \current_shift_inst.control_input_1_cry_6\,
            clk => \N__50187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_7_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46834\,
            in2 => \_gnd_net_\,
            in3 => \N__34162\,
            lcout => \current_shift_inst.control_inputZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_6\,
            carryout => \current_shift_inst.control_input_1_cry_7\,
            clk => \N__50187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_8_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34159\,
            in2 => \_gnd_net_\,
            in3 => \N__34144\,
            lcout => \current_shift_inst.control_inputZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.control_input_1_cry_8\,
            clk => \N__50181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_9_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34141\,
            in2 => \_gnd_net_\,
            in3 => \N__34120\,
            lcout => \current_shift_inst.control_inputZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_8\,
            carryout => \current_shift_inst.control_input_1_cry_9\,
            clk => \N__50181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_10_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34117\,
            in2 => \_gnd_net_\,
            in3 => \N__34099\,
            lcout => \current_shift_inst.control_inputZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_9\,
            carryout => \current_shift_inst.control_input_1_cry_10\,
            clk => \N__50181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_11_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34096\,
            in2 => \_gnd_net_\,
            in3 => \N__34081\,
            lcout => \current_shift_inst.control_inputZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_10\,
            carryout => \current_shift_inst.control_input_1_cry_11\,
            clk => \N__50181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_12_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34078\,
            in2 => \_gnd_net_\,
            in3 => \N__34063\,
            lcout => \current_shift_inst.control_inputZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_11\,
            carryout => \current_shift_inst.control_input_1_cry_12\,
            clk => \N__50181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_13_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34324\,
            in2 => \_gnd_net_\,
            in3 => \N__34306\,
            lcout => \current_shift_inst.control_inputZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_12\,
            carryout => \current_shift_inst.control_input_1_cry_13\,
            clk => \N__50181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_14_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34303\,
            in2 => \_gnd_net_\,
            in3 => \N__34288\,
            lcout => \current_shift_inst.control_inputZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_13\,
            carryout => \current_shift_inst.control_input_1_cry_14\,
            clk => \N__50181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_15_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34285\,
            in2 => \_gnd_net_\,
            in3 => \N__34270\,
            lcout => \current_shift_inst.control_inputZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_14\,
            carryout => \current_shift_inst.control_input_1_cry_15\,
            clk => \N__50181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_16_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34573\,
            in2 => \_gnd_net_\,
            in3 => \N__34258\,
            lcout => \current_shift_inst.control_inputZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.control_input_1_cry_16\,
            clk => \N__50176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_17_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34255\,
            in2 => \_gnd_net_\,
            in3 => \N__34237\,
            lcout => \current_shift_inst.control_inputZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_16\,
            carryout => \current_shift_inst.control_input_1_cry_17\,
            clk => \N__50176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_18_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34492\,
            in2 => \_gnd_net_\,
            in3 => \N__34225\,
            lcout => \current_shift_inst.control_inputZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_17\,
            carryout => \current_shift_inst.control_input_1_cry_18\,
            clk => \N__50176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_19_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34633\,
            in2 => \_gnd_net_\,
            in3 => \N__34213\,
            lcout => \current_shift_inst.control_inputZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_18\,
            carryout => \current_shift_inst.control_input_1_cry_19\,
            clk => \N__50176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_20_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34471\,
            in2 => \_gnd_net_\,
            in3 => \N__34201\,
            lcout => \current_shift_inst.control_inputZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_19\,
            carryout => \current_shift_inst.control_input_1_cry_20\,
            clk => \N__50176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_21_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34522\,
            in2 => \_gnd_net_\,
            in3 => \N__34447\,
            lcout => \current_shift_inst.control_inputZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_20\,
            carryout => \current_shift_inst.control_input_1_cry_21\,
            clk => \N__50176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_22_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34363\,
            in2 => \_gnd_net_\,
            in3 => \N__34432\,
            lcout => \current_shift_inst.control_inputZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_21\,
            carryout => \current_shift_inst.control_input_1_cry_22\,
            clk => \N__50176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_23_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34555\,
            in2 => \_gnd_net_\,
            in3 => \N__34420\,
            lcout => \current_shift_inst.control_inputZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_22\,
            carryout => \current_shift_inst.control_input_1_cry_23\,
            clk => \N__50176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_24_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34618\,
            in2 => \_gnd_net_\,
            in3 => \N__34405\,
            lcout => \current_shift_inst.control_inputZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \current_shift_inst.control_input_1_cry_24\,
            clk => \N__50171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_25_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34402\,
            in2 => \_gnd_net_\,
            in3 => \N__34390\,
            lcout => \current_shift_inst.control_inputZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100110101"
        )
    port map (
            in0 => \N__38629\,
            in1 => \N__34372\,
            in2 => \N__46930\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46901\,
            lcout => \current_shift_inst.N_1355_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101010011"
        )
    port map (
            in0 => \N__34339\,
            in1 => \N__38470\,
            in2 => \N__46929\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__34582\,
            in1 => \N__38716\,
            in2 => \_gnd_net_\,
            in3 => \N__46902\,
            lcout => \current_shift_inst.control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34567\,
            in2 => \N__46931\,
            in3 => \N__39097\,
            lcout => \current_shift_inst.control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38461\,
            in1 => \N__34549\,
            in2 => \_gnd_net_\,
            in3 => \N__46897\,
            lcout => \current_shift_inst.control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__46927\,
            in1 => \_gnd_net_\,
            in2 => \N__38644\,
            in3 => \N__34531\,
            lcout => \current_shift_inst.control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__46771\,
            in1 => \N__46232\,
            in2 => \N__47635\,
            in3 => \N__42907\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46231\,
            in1 => \N__46772\,
            in2 => \N__48064\,
            in3 => \N__45442\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38683\,
            in1 => \N__34498\,
            in2 => \_gnd_net_\,
            in3 => \N__46924\,
            lcout => \current_shift_inst.control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__46233\,
            in1 => \N__46773\,
            in2 => \N__47953\,
            in3 => \N__43089\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__34477\,
            in1 => \N__38656\,
            in2 => \_gnd_net_\,
            in3 => \N__46926\,
            lcout => \current_shift_inst.control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__46925\,
            in1 => \N__34639\,
            in2 => \_gnd_net_\,
            in3 => \N__38668\,
            lcout => \current_shift_inst.control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__34624\,
            in1 => \N__39082\,
            in2 => \_gnd_net_\,
            in3 => \N__46928\,
            lcout => \current_shift_inst.control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46740\,
            in1 => \N__48343\,
            in2 => \N__46342\,
            in3 => \N__43252\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46741\,
            in1 => \N__48427\,
            in2 => \N__46344\,
            in3 => \N__43288\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46739\,
            in1 => \N__48497\,
            in2 => \N__46343\,
            in3 => \N__43024\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34823\,
            in1 => \N__38897\,
            in2 => \_gnd_net_\,
            in3 => \N__34594\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__50158\,
            ce => \N__34726\,
            sr => \N__49691\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34818\,
            in1 => \N__38852\,
            in2 => \_gnd_net_\,
            in3 => \N__34591\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__50158\,
            ce => \N__34726\,
            sr => \N__49691\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34824\,
            in1 => \N__35162\,
            in2 => \_gnd_net_\,
            in3 => \N__34588\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__50158\,
            ce => \N__34726\,
            sr => \N__49691\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34819\,
            in1 => \N__35114\,
            in2 => \_gnd_net_\,
            in3 => \N__34585\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__50158\,
            ce => \N__34726\,
            sr => \N__49691\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34825\,
            in1 => \N__35058\,
            in2 => \_gnd_net_\,
            in3 => \N__34666\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__50158\,
            ce => \N__34726\,
            sr => \N__49691\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34820\,
            in1 => \N__35003\,
            in2 => \_gnd_net_\,
            in3 => \N__34663\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__50158\,
            ce => \N__34726\,
            sr => \N__49691\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34822\,
            in1 => \N__34938\,
            in2 => \_gnd_net_\,
            in3 => \N__34660\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__50158\,
            ce => \N__34726\,
            sr => \N__49691\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34821\,
            in1 => \N__35592\,
            in2 => \_gnd_net_\,
            in3 => \N__34657\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__50158\,
            ce => \N__34726\,
            sr => \N__49691\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34852\,
            in1 => \N__35540\,
            in2 => \_gnd_net_\,
            in3 => \N__34654\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__50154\,
            ce => \N__34739\,
            sr => \N__49700\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34870\,
            in1 => \N__35483\,
            in2 => \_gnd_net_\,
            in3 => \N__34651\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__50154\,
            ce => \N__34739\,
            sr => \N__49700\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34849\,
            in1 => \N__35432\,
            in2 => \_gnd_net_\,
            in3 => \N__34648\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__50154\,
            ce => \N__34739\,
            sr => \N__49700\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34867\,
            in1 => \N__35375\,
            in2 => \_gnd_net_\,
            in3 => \N__34645\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__50154\,
            ce => \N__34739\,
            sr => \N__49700\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34850\,
            in1 => \N__35313\,
            in2 => \_gnd_net_\,
            in3 => \N__34642\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__50154\,
            ce => \N__34739\,
            sr => \N__49700\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34868\,
            in1 => \N__35261\,
            in2 => \_gnd_net_\,
            in3 => \N__34693\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__50154\,
            ce => \N__34739\,
            sr => \N__49700\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34851\,
            in1 => \N__35235\,
            in2 => \_gnd_net_\,
            in3 => \N__34690\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__50154\,
            ce => \N__34739\,
            sr => \N__49700\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34869\,
            in1 => \N__35877\,
            in2 => \_gnd_net_\,
            in3 => \N__34687\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__50154\,
            ce => \N__34739\,
            sr => \N__49700\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34863\,
            in1 => \N__35846\,
            in2 => \_gnd_net_\,
            in3 => \N__34684\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__50150\,
            ce => \N__34741\,
            sr => \N__49704\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34853\,
            in1 => \N__35813\,
            in2 => \_gnd_net_\,
            in3 => \N__34681\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__50150\,
            ce => \N__34741\,
            sr => \N__49704\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34864\,
            in1 => \N__35774\,
            in2 => \_gnd_net_\,
            in3 => \N__34678\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__50150\,
            ce => \N__34741\,
            sr => \N__49704\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34854\,
            in1 => \N__35738\,
            in2 => \_gnd_net_\,
            in3 => \N__34675\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__50150\,
            ce => \N__34741\,
            sr => \N__49704\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34865\,
            in1 => \N__35694\,
            in2 => \_gnd_net_\,
            in3 => \N__34672\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__50150\,
            ce => \N__34741\,
            sr => \N__49704\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34855\,
            in1 => \N__35663\,
            in2 => \_gnd_net_\,
            in3 => \N__34669\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__50150\,
            ce => \N__34741\,
            sr => \N__49704\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34866\,
            in1 => \N__35631\,
            in2 => \_gnd_net_\,
            in3 => \N__34891\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__50150\,
            ce => \N__34741\,
            sr => \N__49704\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34856\,
            in1 => \N__36126\,
            in2 => \_gnd_net_\,
            in3 => \N__34888\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__50150\,
            ce => \N__34741\,
            sr => \N__49704\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34857\,
            in1 => \N__36089\,
            in2 => \_gnd_net_\,
            in3 => \N__34885\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__50145\,
            ce => \N__34740\,
            sr => \N__49709\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34861\,
            in1 => \N__36050\,
            in2 => \_gnd_net_\,
            in3 => \N__34882\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__50145\,
            ce => \N__34740\,
            sr => \N__49709\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34858\,
            in1 => \N__36020\,
            in2 => \_gnd_net_\,
            in3 => \N__34879\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__50145\,
            ce => \N__34740\,
            sr => \N__49709\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34862\,
            in1 => \N__35966\,
            in2 => \_gnd_net_\,
            in3 => \N__34876\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__50145\,
            ce => \N__34740\,
            sr => \N__49709\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34859\,
            in1 => \N__35994\,
            in2 => \_gnd_net_\,
            in3 => \N__34873\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__50145\,
            ce => \N__34740\,
            sr => \N__49709\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__35943\,
            in1 => \N__34860\,
            in2 => \_gnd_net_\,
            in3 => \N__34744\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50145\,
            ce => \N__34740\,
            sr => \N__49709\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__35564\,
            in1 => \N__35202\,
            in2 => \N__38962\,
            in3 => \N__38831\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRMG72_7_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34972\,
            in2 => \N__35218\,
            in3 => \N__35040\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38904\,
            in2 => \N__35167\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__50137\,
            ce => \N__38811\,
            sr => \N__49726\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38859\,
            in2 => \N__35119\,
            in3 => \N__35170\,
            lcout => \delay_measurement_inst.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__50137\,
            ce => \N__38811\,
            sr => \N__49726\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35166\,
            in2 => \N__35070\,
            in3 => \N__35122\,
            lcout => \delay_measurement_inst.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__50137\,
            ce => \N__38811\,
            sr => \N__49726\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35118\,
            in2 => \N__35014\,
            in3 => \N__35074\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__50137\,
            ce => \N__38811\,
            sr => \N__49726\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34944\,
            in2 => \N__35071\,
            in3 => \N__35017\,
            lcout => \delay_measurement_inst.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__50137\,
            ce => \N__38811\,
            sr => \N__49726\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35013\,
            in2 => \N__35604\,
            in3 => \N__34948\,
            lcout => \delay_measurement_inst.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__50137\,
            ce => \N__38811\,
            sr => \N__49726\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34945\,
            in2 => \N__35545\,
            in3 => \N__34894\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__50137\,
            ce => \N__38811\,
            sr => \N__49726\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35490\,
            in2 => \N__35605\,
            in3 => \N__35548\,
            lcout => \delay_measurement_inst.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__50137\,
            ce => \N__38811\,
            sr => \N__49726\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35544\,
            in2 => \N__35437\,
            in3 => \N__35497\,
            lcout => \delay_measurement_inst.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_14_27_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__50134\,
            ce => \N__38810\,
            sr => \N__49731\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35494\,
            in2 => \N__35380\,
            in3 => \N__35440\,
            lcout => \delay_measurement_inst.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__50134\,
            ce => \N__38810\,
            sr => \N__49731\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35436\,
            in2 => \N__35325\,
            in3 => \N__35383\,
            lcout => \delay_measurement_inst.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__50134\,
            ce => \N__38810\,
            sr => \N__49731\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35379\,
            in2 => \N__35268\,
            in3 => \N__35329\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__50134\,
            ce => \N__38810\,
            sr => \N__49731\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35241\,
            in2 => \N__35326\,
            in3 => \N__35272\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__50134\,
            ce => \N__38810\,
            sr => \N__49731\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35883\,
            in2 => \N__35269\,
            in3 => \N__35245\,
            lcout => \delay_measurement_inst.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__50134\,
            ce => \N__38810\,
            sr => \N__49731\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35242\,
            in2 => \N__35859\,
            in3 => \N__35221\,
            lcout => \delay_measurement_inst.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__50134\,
            ce => \N__38810\,
            sr => \N__49731\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35884\,
            in2 => \N__35826\,
            in3 => \N__35863\,
            lcout => \delay_measurement_inst.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__50134\,
            ce => \N__38810\,
            sr => \N__49731\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35860\,
            in2 => \N__35779\,
            in3 => \N__35830\,
            lcout => \delay_measurement_inst.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_14_28_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__50132\,
            ce => \N__38809\,
            sr => \N__49736\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35827\,
            in2 => \N__35743\,
            in3 => \N__35782\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__50132\,
            ce => \N__38809\,
            sr => \N__49736\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35778\,
            in2 => \N__35706\,
            in3 => \N__35746\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__50132\,
            ce => \N__38809\,
            sr => \N__49736\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35742\,
            in2 => \N__35670\,
            in3 => \N__35710\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__50132\,
            ce => \N__38809\,
            sr => \N__49736\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35637\,
            in2 => \N__35707\,
            in3 => \N__35674\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__50132\,
            ce => \N__38809\,
            sr => \N__49736\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36132\,
            in2 => \N__35671\,
            in3 => \N__35641\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__50132\,
            ce => \N__38809\,
            sr => \N__49736\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35638\,
            in2 => \N__36100\,
            in3 => \N__35608\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__50132\,
            ce => \N__38809\,
            sr => \N__49736\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36133\,
            in2 => \N__36063\,
            in3 => \N__36103\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__50132\,
            ce => \N__38809\,
            sr => \N__49736\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_14_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36099\,
            in2 => \N__36025\,
            in3 => \N__36067\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_14_29_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__50130\,
            ce => \N__38808\,
            sr => \N__49738\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36064\,
            in2 => \N__35971\,
            in3 => \N__36028\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__50130\,
            ce => \N__38808\,
            sr => \N__49738\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36024\,
            in2 => \N__36001\,
            in3 => \N__35974\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__50130\,
            ce => \N__38808\,
            sr => \N__49738\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35970\,
            in2 => \N__35947\,
            in3 => \N__35920\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__50130\,
            ce => \N__38808\,
            sr => \N__49738\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35917\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50130\,
            ce => \N__38808\,
            sr => \N__49738\
        );

    \SB_DFF_inst_DELAY_TR1_LC_15_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35899\,
            lcout => delay_tr_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR2_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35890\,
            lcout => delay_tr_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_15_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__39187\,
            in1 => \N__39208\,
            in2 => \N__49791\,
            in3 => \N__39169\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_0_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__39188\,
            in1 => \N__39206\,
            in2 => \_gnd_net_\,
            in3 => \N__39168\,
            lcout => \delay_measurement_inst.tr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50267\,
            ce => \N__36415\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNITAU01_13_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44079\,
            in1 => \N__36322\,
            in2 => \N__43588\,
            in3 => \N__36286\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNITAU01Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000111"
        )
    port map (
            in0 => \N__39505\,
            in1 => \N__45124\,
            in2 => \N__44933\,
            in3 => \N__45338\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50252\,
            ce => 'H',
            sr => \N__49612\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIC46U_6_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44051\,
            in1 => \N__36276\,
            in2 => \N__39392\,
            in3 => \N__36247\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIC46UZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI8V4U_5_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44050\,
            in1 => \N__36240\,
            in2 => \N__36532\,
            in3 => \N__36211\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI8V4UZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI4Q3U_4_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44049\,
            in1 => \N__36204\,
            in2 => \N__39286\,
            in3 => \N__36175\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI4Q3UZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43569\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIKE8U_8_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44053\,
            in1 => \N__36168\,
            in2 => \N__39361\,
            in3 => \N__36139\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIKE8UZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43528\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIG97U_7_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44052\,
            in1 => \N__36682\,
            in2 => \N__40881\,
            in3 => \N__36655\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIG97UZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIOJ9U_9_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__43468\,
            in1 => \N__44054\,
            in2 => \N__36649\,
            in3 => \N__36616\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIOJ9UZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIA1B41_10_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44055\,
            in1 => \N__36609\,
            in2 => \N__43536\,
            in3 => \N__36580\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIA1B41Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIP5T01_12_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__43625\,
            in1 => \N__44056\,
            in2 => \N__36574\,
            in3 => \N__36538\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIP5T01Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41718\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36531\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIL0S01_11_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__36486\,
            in1 => \N__43983\,
            in2 => \N__44203\,
            in3 => \N__36457\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIL0S01Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIDGBQ_22_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43987\,
            in1 => \N__36450\,
            in2 => \N__40207\,
            in3 => \N__36421\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIDGBQZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIGNK3_0_26_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43982\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIS2EP_19_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43986\,
            in1 => \N__36952\,
            in2 => \N__36928\,
            in3 => \N__36877\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIS2EPZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNICE9P_15_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__41728\,
            in1 => \N__43984\,
            in2 => \N__36871\,
            in3 => \N__36861\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNICE9PZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36827\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37115\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIGJAP_16_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__43985\,
            in1 => \N__36778\,
            in2 => \N__41674\,
            in3 => \N__36771\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIGJAPZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIHLCQ_23_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44068\,
            in1 => \N__36738\,
            in2 => \N__40150\,
            in3 => \N__36709\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIHLCQZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__36703\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44066\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8J_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__44070\,
            in1 => \N__44453\,
            in2 => \N__36691\,
            in3 => \N__36688\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJ_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__37234\,
            in1 => \N__44073\,
            in2 => \N__44651\,
            in3 => \N__37210\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7J_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__44069\,
            in1 => \N__37204\,
            in2 => \N__39492\,
            in3 => \N__37180\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJ_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101101111011"
        )
    port map (
            in0 => \N__37173\,
            in1 => \N__44072\,
            in2 => \N__37156\,
            in3 => \N__41338\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIENGP_20_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44067\,
            in1 => \N__37146\,
            in2 => \N__37120\,
            in3 => \N__37075\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIENGPZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9J_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__37069\,
            in1 => \N__44071\,
            in2 => \N__44581\,
            in3 => \N__37045\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50328\,
            in2 => \N__41610\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__50222\,
            ce => \N__49811\,
            sr => \N__49625\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44332\,
            in2 => \N__42090\,
            in3 => \N__36976\,
            lcout => \delay_measurement_inst.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__50222\,
            ce => \N__49811\,
            sr => \N__49625\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42063\,
            in2 => \N__41611\,
            in3 => \N__36955\,
            lcout => \delay_measurement_inst.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__50222\,
            ce => \N__49811\,
            sr => \N__49625\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42042\,
            in2 => \N__42091\,
            in3 => \N__37435\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__50222\,
            ce => \N__49811\,
            sr => \N__49625\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42064\,
            in2 => \N__42018\,
            in3 => \N__37408\,
            lcout => \delay_measurement_inst.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__50222\,
            ce => \N__49811\,
            sr => \N__49625\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42043\,
            in2 => \N__41991\,
            in3 => \N__37384\,
            lcout => \delay_measurement_inst.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__50222\,
            ce => \N__49811\,
            sr => \N__49625\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41965\,
            in2 => \N__42019\,
            in3 => \N__37330\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__50222\,
            ce => \N__49811\,
            sr => \N__49625\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41938\,
            in2 => \N__41992\,
            in3 => \N__37306\,
            lcout => \delay_measurement_inst.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__50222\,
            ce => \N__49811\,
            sr => \N__49625\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41964\,
            in2 => \N__41907\,
            in3 => \N__37285\,
            lcout => \delay_measurement_inst.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__50212\,
            ce => \N__49812\,
            sr => \N__49630\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41937\,
            in2 => \N__41880\,
            in3 => \N__37261\,
            lcout => \delay_measurement_inst.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__50212\,
            ce => \N__49812\,
            sr => \N__49630\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42300\,
            in2 => \N__41908\,
            in3 => \N__37237\,
            lcout => \delay_measurement_inst.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__50212\,
            ce => \N__49812\,
            sr => \N__49630\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42276\,
            in2 => \N__41881\,
            in3 => \N__37702\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__50212\,
            ce => \N__49812\,
            sr => \N__49630\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42301\,
            in2 => \N__42255\,
            in3 => \N__37654\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__50212\,
            ce => \N__49812\,
            sr => \N__49630\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42277\,
            in2 => \N__42228\,
            in3 => \N__37618\,
            lcout => \delay_measurement_inst.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__50212\,
            ce => \N__49812\,
            sr => \N__49630\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42202\,
            in2 => \N__42256\,
            in3 => \N__37576\,
            lcout => \delay_measurement_inst.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__50212\,
            ce => \N__49812\,
            sr => \N__49630\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42172\,
            in2 => \N__42229\,
            in3 => \N__37537\,
            lcout => \delay_measurement_inst.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__50212\,
            ce => \N__49812\,
            sr => \N__49630\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42201\,
            in2 => \N__42144\,
            in3 => \N__37498\,
            lcout => \delay_measurement_inst.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__50208\,
            ce => \N__49813\,
            sr => \N__49639\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42171\,
            in2 => \N__42117\,
            in3 => \N__37495\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__50208\,
            ce => \N__49813\,
            sr => \N__49639\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42525\,
            in2 => \N__42145\,
            in3 => \N__37492\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__50208\,
            ce => \N__49813\,
            sr => \N__49639\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42504\,
            in2 => \N__42118\,
            in3 => \N__37489\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__50208\,
            ce => \N__49813\,
            sr => \N__49639\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42526\,
            in2 => \N__42483\,
            in3 => \N__37822\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__50208\,
            ce => \N__49813\,
            sr => \N__49639\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42505\,
            in2 => \N__42456\,
            in3 => \N__37813\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__50208\,
            ce => \N__49813\,
            sr => \N__49639\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42430\,
            in2 => \N__42484\,
            in3 => \N__37804\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__50208\,
            ce => \N__49813\,
            sr => \N__49639\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42403\,
            in2 => \N__42457\,
            in3 => \N__37795\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__50208\,
            ce => \N__49813\,
            sr => \N__49639\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42429\,
            in2 => \N__42372\,
            in3 => \N__37783\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__50202\,
            ce => \N__49814\,
            sr => \N__49645\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42402\,
            in2 => \N__42345\,
            in3 => \N__37771\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__50202\,
            ce => \N__49814\,
            sr => \N__49645\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42319\,
            in2 => \N__42373\,
            in3 => \N__37759\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__50202\,
            ce => \N__49814\,
            sr => \N__49645\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42655\,
            in2 => \N__42346\,
            in3 => \N__37741\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__50202\,
            ce => \N__49814\,
            sr => \N__49645\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37939\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50202\,
            ce => \N__49814\,
            sr => \N__49645\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45360\,
            in2 => \N__37852\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40357\,
            in2 => \N__38380\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47125\,
            in2 => \N__38384\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40465\,
            in2 => \N__38381\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38326\,
            in2 => \N__40447\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40453\,
            in2 => \N__38382\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45469\,
            in2 => \N__38385\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40459\,
            in2 => \N__38383\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40525\,
            in2 => \N__38375\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40489\,
            in2 => \N__38379\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40495\,
            in2 => \N__38372\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40507\,
            in2 => \N__38376\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40519\,
            in2 => \N__38373\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40531\,
            in2 => \N__38377\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40501\,
            in2 => \N__38374\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40513\,
            in2 => \N__38378\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40609\,
            in2 => \N__38289\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40603\,
            in2 => \N__38293\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45409\,
            in2 => \N__38290\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40483\,
            in2 => \N__38294\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40654\,
            in2 => \N__38291\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38200\,
            in2 => \N__40648\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40597\,
            in2 => \N__38292\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40567\,
            in2 => \N__38295\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40552\,
            in2 => \N__38280\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40666\,
            in2 => \N__38284\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40540\,
            in2 => \N__38281\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40546\,
            in2 => \N__38285\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40615\,
            in2 => \N__38282\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40729\,
            in2 => \N__38286\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43186\,
            in2 => \N__38283\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46749\,
            in2 => \_gnd_net_\,
            in3 => \N__37996\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37993\,
            in2 => \N__37974\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40387\,
            in2 => \N__40425\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37951\,
            in2 => \N__46255\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40477\,
            in2 => \N__46258\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40717\,
            in2 => \N__46256\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40660\,
            in2 => \N__46259\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47062\,
            in2 => \N__46257\,
            in3 => \N__38464\,
            lcout => \current_shift_inst.un38_control_input_0_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47383\,
            in2 => \N__46260\,
            in3 => \N__38452\,
            lcout => \current_shift_inst.un38_control_input_0_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40627\,
            in2 => \N__46325\,
            in3 => \N__38437\,
            lcout => \current_shift_inst.un38_control_input_0_s1_8\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40579\,
            in2 => \N__46329\,
            in3 => \N__38422\,
            lcout => \current_shift_inst.un38_control_input_0_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40735\,
            in2 => \N__46326\,
            in3 => \N__38404\,
            lcout => \current_shift_inst.un38_control_input_0_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40723\,
            in2 => \N__46330\,
            in3 => \N__38401\,
            lcout => \current_shift_inst.un38_control_input_0_s1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40561\,
            in2 => \N__46327\,
            in3 => \N__38599\,
            lcout => \current_shift_inst.un38_control_input_0_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40621\,
            in2 => \N__46331\,
            in3 => \N__38596\,
            lcout => \current_shift_inst.un38_control_input_0_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40687\,
            in2 => \N__46328\,
            in3 => \N__38578\,
            lcout => \current_shift_inst.un38_control_input_0_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40753\,
            in2 => \N__46332\,
            in3 => \N__38560\,
            lcout => \current_shift_inst.un38_control_input_0_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41263\,
            in2 => \N__46366\,
            in3 => \N__38542\,
            lcout => \current_shift_inst.un38_control_input_0_s1_16\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40699\,
            in2 => \N__46273\,
            in3 => \N__38524\,
            lcout => \current_shift_inst.un38_control_input_0_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40813\,
            in2 => \N__46367\,
            in3 => \N__38506\,
            lcout => \current_shift_inst.un38_control_input_0_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40693\,
            in2 => \N__46274\,
            in3 => \N__38488\,
            lcout => \current_shift_inst.un38_control_input_0_s1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40801\,
            in2 => \N__46368\,
            in3 => \N__38737\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41275\,
            in2 => \N__46275\,
            in3 => \N__38719\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40795\,
            in2 => \N__46369\,
            in3 => \N__38704\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40807\,
            in2 => \N__46276\,
            in3 => \N__38686\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40639\,
            in2 => \N__46375\,
            in3 => \N__38671\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40759\,
            in2 => \N__46370\,
            in3 => \N__38659\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40765\,
            in2 => \N__46376\,
            in3 => \N__38647\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41269\,
            in2 => \N__46371\,
            in3 => \N__38632\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46283\,
            in2 => \N__40747\,
            in3 => \N__38617\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40789\,
            in2 => \N__46372\,
            in3 => \N__39085\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40776\,
            in2 => \N__46377\,
            in3 => \N__39070\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_2_25_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__46800\,
            in1 => \N__46315\,
            in2 => \_gnd_net_\,
            in3 => \N__39067\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39048\,
            in1 => \N__39018\,
            in2 => \N__38991\,
            in3 => \N__38961\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38911\,
            lcout => \delay_measurement_inst.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50140\,
            ce => \N__38812\,
            sr => \N__49717\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38863\,
            lcout => \delay_measurement_inst.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50140\,
            ce => \N__38812\,
            sr => \N__49717\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_1_3_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41244\,
            in2 => \_gnd_net_\,
            in3 => \N__41256\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_1_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40902\,
            in1 => \N__41232\,
            in2 => \N__38791\,
            in3 => \N__38788\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_16_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39134\,
            in2 => \_gnd_net_\,
            in3 => \N__39115\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_304_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_16_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__39189\,
            in1 => \N__39207\,
            in2 => \_gnd_net_\,
            in3 => \N__39167\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => 'H',
            sr => \N__49603\
        );

    \delay_measurement_inst.prev_tr_sig_LC_16_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39190\,
            lcout => \delay_measurement_inst.prev_tr_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => 'H',
            sr => \N__49603\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_16_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__39151\,
            in1 => \N__39138\,
            in2 => \_gnd_net_\,
            in3 => \N__39118\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => 'H',
            sr => \N__49603\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39116\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__39150\,
            in1 => \N__39139\,
            in2 => \_gnd_net_\,
            in3 => \N__39117\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_305_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__45112\,
            in1 => \N__45340\,
            in2 => \_gnd_net_\,
            in3 => \N__39268\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50263\,
            ce => 'H',
            sr => \N__49608\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45136\,
            in1 => \N__45303\,
            in2 => \N__44935\,
            in3 => \N__39613\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49609\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__45301\,
            in1 => \N__45137\,
            in2 => \_gnd_net_\,
            in3 => \N__39658\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49609\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45135\,
            in1 => \N__45302\,
            in2 => \N__44934\,
            in3 => \N__39862\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50257\,
            ce => 'H',
            sr => \N__49609\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39425\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40854\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39377\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39331\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41428\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39309\,
            in2 => \N__39310\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39292\,
            in2 => \N__39285\,
            in3 => \N__39259\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39256\,
            in2 => \N__39250\,
            in3 => \N__39226\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39673\,
            in2 => \N__39667\,
            in3 => \N__39649\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39646\,
            in2 => \N__39640\,
            in3 => \N__39631\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39628\,
            in2 => \N__39622\,
            in3 => \N__39604\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39601\,
            in2 => \N__39595\,
            in3 => \N__39580\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39577\,
            in2 => \N__39571\,
            in3 => \N__39553\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39550\,
            in2 => \N__44152\,
            in3 => \N__39541\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39538\,
            in2 => \N__41473\,
            in3 => \N__39532\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39529\,
            in2 => \N__39517\,
            in3 => \N__39496\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43825\,
            in2 => \N__44218\,
            in3 => \N__39814\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39811\,
            in2 => \N__39805\,
            in3 => \N__39796\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39793\,
            in2 => \N__41629\,
            in3 => \N__39787\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44227\,
            in2 => \N__44095\,
            in3 => \N__39772\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41530\,
            in2 => \N__41482\,
            in3 => \N__39757\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39754\,
            in2 => \N__39748\,
            in3 => \N__39724\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39721\,
            in2 => \N__39715\,
            in3 => \N__39694\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41812\,
            in2 => \N__39691\,
            in3 => \N__39676\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39925\,
            in2 => \N__40351\,
            in3 => \N__39919\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40339\,
            in2 => \N__39916\,
            in3 => \N__39907\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40288\,
            in2 => \N__39952\,
            in3 => \N__39904\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41398\,
            in2 => \N__39901\,
            in3 => \N__39886\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39883\,
            in2 => \N__39877\,
            in3 => \N__39853\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39850\,
            in2 => \N__44407\,
            in3 => \N__39844\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39841\,
            in2 => \N__44533\,
            in3 => \N__39826\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39823\,
            in2 => \N__40828\,
            in3 => \N__39817\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40087\,
            in2 => \N__44593\,
            in3 => \N__40081\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40078\,
            in2 => \N__40066\,
            in3 => \N__40045\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39935\,
            in2 => \N__44473\,
            in3 => \N__40042\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39958\,
            in2 => \N__39940\,
            in3 => \N__40030\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39939\,
            in2 => \N__40027\,
            in3 => \N__40003\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43998\,
            in1 => \N__44852\,
            in2 => \_gnd_net_\,
            in3 => \N__40000\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39997\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40240\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIGNK3_26_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43997\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40182\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40117\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNICIEQ_24_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43996\,
            in1 => \N__40326\,
            in2 => \N__40258\,
            in3 => \N__40300\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNICIEQZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011111110"
        )
    port map (
            in0 => \N__45249\,
            in1 => \N__45132\,
            in2 => \N__44923\,
            in3 => \N__40279\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49631\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45130\,
            in1 => \N__45250\,
            in2 => \N__44911\,
            in3 => \N__40216\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49631\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45131\,
            in1 => \N__45251\,
            in2 => \N__44912\,
            in3 => \N__40159\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50213\,
            ce => 'H',
            sr => \N__49631\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40372\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46682\,
            in1 => \N__47478\,
            in2 => \N__46374\,
            in3 => \N__42576\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__42577\,
            in1 => \N__46681\,
            in2 => \N__47482\,
            in3 => \N__46301\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47223\,
            in1 => \N__47477\,
            in2 => \_gnd_net_\,
            in3 => \N__42575\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47226\,
            in1 => \N__47829\,
            in2 => \_gnd_net_\,
            in3 => \N__47399\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47224\,
            in1 => \N__47901\,
            in2 => \_gnd_net_\,
            in3 => \N__42551\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47225\,
            in1 => \N__47449\,
            in2 => \_gnd_net_\,
            in3 => \N__45563\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__46679\,
            in1 => \N__42591\,
            in2 => \N__40426\,
            in3 => \N__40374\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48778\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50203\,
            ce => \N__48267\,
            sr => \N__49646\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__40375\,
            in1 => \N__46678\,
            in2 => \N__42595\,
            in3 => \N__40424\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__47265\,
            in1 => \N__42590\,
            in2 => \_gnd_net_\,
            in3 => \N__40373\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__43280\,
            in1 => \N__46680\,
            in2 => \_gnd_net_\,
            in3 => \N__48426\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47586\,
            in1 => \N__47280\,
            in2 => \_gnd_net_\,
            in3 => \N__42869\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47277\,
            in1 => \N__47795\,
            in2 => \_gnd_net_\,
            in3 => \N__42986\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47630\,
            in1 => \N__47279\,
            in2 => \_gnd_net_\,
            in3 => \N__42899\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47281\,
            in1 => \N__48188\,
            in2 => \_gnd_net_\,
            in3 => \N__42806\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47267\,
            in1 => \N__47673\,
            in2 => \_gnd_net_\,
            in3 => \N__47111\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48233\,
            in1 => \N__47268\,
            in2 => \_gnd_net_\,
            in3 => \N__42839\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47266\,
            in1 => \N__47709\,
            in2 => \_gnd_net_\,
            in3 => \N__42929\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47278\,
            in1 => \N__47750\,
            in2 => \_gnd_net_\,
            in3 => \N__42959\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47273\,
            in1 => \N__48018\,
            in2 => \_gnd_net_\,
            in3 => \N__43127\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47269\,
            in1 => \N__48144\,
            in2 => \_gnd_net_\,
            in3 => \N__45503\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47272\,
            in1 => \N__48099\,
            in2 => \_gnd_net_\,
            in3 => \N__43364\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47270\,
            in1 => \N__48578\,
            in2 => \_gnd_net_\,
            in3 => \N__43041\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46704\,
            in1 => \N__48019\,
            in2 => \N__46324\,
            in3 => \N__43128\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__46702\,
            in1 => \N__42960\,
            in2 => \N__46229\,
            in3 => \N__47751\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48537\,
            in1 => \N__47271\,
            in2 => \_gnd_net_\,
            in3 => \N__43163\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46703\,
            in1 => \N__47631\,
            in2 => \N__46230\,
            in3 => \N__42900\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47275\,
            in1 => \N__48498\,
            in2 => \_gnd_net_\,
            in3 => \N__43016\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46690\,
            in1 => \N__48381\,
            in2 => \_gnd_net_\,
            in3 => \N__43313\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__43107\,
            in1 => \N__46691\,
            in2 => \N__47986\,
            in3 => \N__46152\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46689\,
            in1 => \N__48465\,
            in2 => \_gnd_net_\,
            in3 => \N__43694\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__42559\,
            in1 => \N__46688\,
            in2 => \N__46290\,
            in3 => \N__47900\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47276\,
            in1 => \N__47981\,
            in2 => \_gnd_net_\,
            in3 => \N__43106\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47274\,
            in1 => \N__47952\,
            in2 => \_gnd_net_\,
            in3 => \N__43076\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__43017\,
            in1 => \N__46799\,
            in2 => \N__48502\,
            in3 => \N__46098\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46692\,
            in1 => \N__47796\,
            in2 => \N__46293\,
            in3 => \N__43000\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46687\,
            in1 => \N__47585\,
            in2 => \N__46320\,
            in3 => \N__42876\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48341\,
            in1 => \N__46684\,
            in2 => \_gnd_net_\,
            in3 => \N__43241\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__43242\,
            in1 => \N__46694\,
            in2 => \N__46319\,
            in3 => \N__48342\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46693\,
            in1 => \N__47708\,
            in2 => \N__46291\,
            in3 => \N__42940\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46685\,
            in1 => \N__48302\,
            in2 => \_gnd_net_\,
            in3 => \N__43217\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__47116\,
            in1 => \N__46686\,
            in2 => \N__46292\,
            in3 => \N__47672\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46683\,
            in1 => \N__47447\,
            in2 => \N__46321\,
            in3 => \N__45574\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46813\,
            in1 => \N__48307\,
            in2 => \N__46296\,
            in3 => \N__43224\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46810\,
            in1 => \N__48100\,
            in2 => \N__46297\,
            in3 => \N__43375\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46701\,
            in1 => \N__48017\,
            in2 => \N__46334\,
            in3 => \N__43132\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46809\,
            in1 => \N__48234\,
            in2 => \N__46294\,
            in3 => \N__42850\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46700\,
            in1 => \N__48056\,
            in2 => \N__46333\,
            in3 => \N__45441\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46812\,
            in1 => \N__48538\,
            in2 => \N__46295\,
            in3 => \N__43171\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47985\,
            in1 => \N__46811\,
            in2 => \N__46335\,
            in3 => \N__43111\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46697\,
            in1 => \N__48579\,
            in2 => \N__46302\,
            in3 => \N__43053\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__43225\,
            in1 => \N__46817\,
            in2 => \N__46303\,
            in3 => \N__48303\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46699\,
            in2 => \_gnd_net_\,
            in3 => \N__43198\,
            lcout => \current_shift_inst.un4_control_input_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46698\,
            in1 => \N__48419\,
            in2 => \N__46305\,
            in3 => \N__43287\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46816\,
            in1 => \N__48466\,
            in2 => \N__46323\,
            in3 => \N__43705\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46695\,
            in1 => \N__48189\,
            in2 => \N__46304\,
            in3 => \N__42820\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47948\,
            in1 => \N__46696\,
            in2 => \N__46322\,
            in3 => \N__43090\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46815\,
            in1 => \N__48382\,
            in2 => \N__46378\,
            in3 => \N__43324\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46814\,
            in1 => \N__48145\,
            in2 => \N__46373\,
            in3 => \N__45517\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_29_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__41187\,
            in1 => \N__41257\,
            in2 => \_gnd_net_\,
            in3 => \N__41050\,
            lcout => measured_delay_hc_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50146\,
            ce => 'H',
            sr => \N__49710\
        );

    \delay_measurement_inst.delay_hc_reg_30_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__41042\,
            in1 => \_gnd_net_\,
            in2 => \N__41221\,
            in3 => \N__41245\,
            lcout => measured_delay_hc_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50141\,
            ce => 'H',
            sr => \N__49718\
        );

    \delay_measurement_inst.delay_hc_reg_27_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__41233\,
            in1 => \N__41214\,
            in2 => \_gnd_net_\,
            in3 => \N__41040\,
            lcout => measured_delay_hc_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50141\,
            ce => 'H',
            sr => \N__49718\
        );

    \delay_measurement_inst.delay_hc_reg_28_LC_16_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__40903\,
            in1 => \N__41215\,
            in2 => \_gnd_net_\,
            in3 => \N__41041\,
            lcout => measured_delay_hc_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50141\,
            ce => 'H',
            sr => \N__49718\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__45138\,
            in1 => \N__45339\,
            in2 => \_gnd_net_\,
            in3 => \N__40891\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50268\,
            ce => 'H',
            sr => \N__49607\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41319\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45134\,
            in1 => \N__45281\,
            in2 => \N__44883\,
            in3 => \N__41584\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50258\,
            ce => 'H',
            sr => \N__49610\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIOTCP_18_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44083\,
            in1 => \N__41571\,
            in2 => \N__41524\,
            in3 => \N__41542\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIOTCPZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41519\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43612\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111110011"
        )
    port map (
            in0 => \N__45133\,
            in1 => \N__44768\,
            in2 => \N__45321\,
            in3 => \N__41464\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50253\,
            ce => 'H',
            sr => \N__49613\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIGNFQ_25_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44082\,
            in1 => \N__41391\,
            in2 => \N__41453\,
            in3 => \N__41410\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIGNFQZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIFMK3_25_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41390\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45046\,
            in1 => \N__45322\,
            in2 => \N__44810\,
            in3 => \N__41353\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50247\,
            ce => 'H',
            sr => \N__49614\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45047\,
            in1 => \N__45323\,
            in2 => \N__44811\,
            in3 => \N__41284\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50247\,
            ce => 'H',
            sr => \N__49614\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI9BAQ_21_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__41854\,
            in1 => \N__44077\,
            in2 => \N__41778\,
            in3 => \N__41841\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI9BAQZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45126\,
            in1 => \N__45305\,
            in2 => \N__44866\,
            in3 => \N__41806\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50241\,
            ce => 'H',
            sr => \N__49617\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45125\,
            in1 => \N__45304\,
            in2 => \N__44865\,
            in3 => \N__41746\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50241\,
            ce => 'H',
            sr => \N__49617\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111011100"
        )
    port map (
            in0 => \N__41680\,
            in1 => \N__44799\,
            in2 => \N__45139\,
            in3 => \N__45306\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50241\,
            ce => 'H',
            sr => \N__49617\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41640\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42780\,
            in1 => \N__50321\,
            in2 => \_gnd_net_\,
            in3 => \N__41617\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__50235\,
            ce => \N__42623\,
            sr => \N__49618\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42776\,
            in1 => \N__44327\,
            in2 => \_gnd_net_\,
            in3 => \N__41614\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__50235\,
            ce => \N__42623\,
            sr => \N__49618\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42781\,
            in1 => \N__41603\,
            in2 => \_gnd_net_\,
            in3 => \N__41587\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__50235\,
            ce => \N__42623\,
            sr => \N__49618\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42777\,
            in1 => \N__42083\,
            in2 => \_gnd_net_\,
            in3 => \N__42067\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__50235\,
            ce => \N__42623\,
            sr => \N__49618\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42782\,
            in1 => \N__42062\,
            in2 => \_gnd_net_\,
            in3 => \N__42046\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__50235\,
            ce => \N__42623\,
            sr => \N__49618\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42778\,
            in1 => \N__42036\,
            in2 => \_gnd_net_\,
            in3 => \N__42022\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__50235\,
            ce => \N__42623\,
            sr => \N__49618\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42783\,
            in1 => \N__42011\,
            in2 => \_gnd_net_\,
            in3 => \N__41995\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__50235\,
            ce => \N__42623\,
            sr => \N__49618\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42779\,
            in1 => \N__41984\,
            in2 => \_gnd_net_\,
            in3 => \N__41968\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__50235\,
            ce => \N__42623\,
            sr => \N__49618\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42775\,
            in1 => \N__41960\,
            in2 => \_gnd_net_\,
            in3 => \N__41941\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__50230\,
            ce => \N__42639\,
            sr => \N__49622\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42771\,
            in1 => \N__41927\,
            in2 => \_gnd_net_\,
            in3 => \N__41911\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__50230\,
            ce => \N__42639\,
            sr => \N__49622\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42772\,
            in1 => \N__41900\,
            in2 => \_gnd_net_\,
            in3 => \N__41884\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__50230\,
            ce => \N__42639\,
            sr => \N__49622\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42768\,
            in1 => \N__41873\,
            in2 => \_gnd_net_\,
            in3 => \N__41857\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__50230\,
            ce => \N__42639\,
            sr => \N__49622\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42773\,
            in1 => \N__42294\,
            in2 => \_gnd_net_\,
            in3 => \N__42280\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__50230\,
            ce => \N__42639\,
            sr => \N__49622\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42769\,
            in1 => \N__42275\,
            in2 => \_gnd_net_\,
            in3 => \N__42259\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__50230\,
            ce => \N__42639\,
            sr => \N__49622\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42774\,
            in1 => \N__42248\,
            in2 => \_gnd_net_\,
            in3 => \N__42232\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__50230\,
            ce => \N__42639\,
            sr => \N__49622\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42770\,
            in1 => \N__42221\,
            in2 => \_gnd_net_\,
            in3 => \N__42205\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__50230\,
            ce => \N__42639\,
            sr => \N__49622\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42764\,
            in1 => \N__42191\,
            in2 => \_gnd_net_\,
            in3 => \N__42175\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__50223\,
            ce => \N__42638\,
            sr => \N__49626\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42784\,
            in1 => \N__42167\,
            in2 => \_gnd_net_\,
            in3 => \N__42148\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__50223\,
            ce => \N__42638\,
            sr => \N__49626\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42765\,
            in1 => \N__42137\,
            in2 => \_gnd_net_\,
            in3 => \N__42121\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__50223\,
            ce => \N__42638\,
            sr => \N__49626\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42785\,
            in1 => \N__42110\,
            in2 => \_gnd_net_\,
            in3 => \N__42094\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__50223\,
            ce => \N__42638\,
            sr => \N__49626\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42766\,
            in1 => \N__42524\,
            in2 => \_gnd_net_\,
            in3 => \N__42508\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__50223\,
            ce => \N__42638\,
            sr => \N__49626\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42786\,
            in1 => \N__42503\,
            in2 => \_gnd_net_\,
            in3 => \N__42487\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__50223\,
            ce => \N__42638\,
            sr => \N__49626\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42767\,
            in1 => \N__42476\,
            in2 => \_gnd_net_\,
            in3 => \N__42460\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__50223\,
            ce => \N__42638\,
            sr => \N__49626\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42787\,
            in1 => \N__42449\,
            in2 => \_gnd_net_\,
            in3 => \N__42433\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__50223\,
            ce => \N__42638\,
            sr => \N__49626\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42758\,
            in1 => \N__42425\,
            in2 => \_gnd_net_\,
            in3 => \N__42406\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__50214\,
            ce => \N__42640\,
            sr => \N__49632\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42762\,
            in1 => \N__42392\,
            in2 => \_gnd_net_\,
            in3 => \N__42376\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__50214\,
            ce => \N__42640\,
            sr => \N__49632\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42759\,
            in1 => \N__42365\,
            in2 => \_gnd_net_\,
            in3 => \N__42349\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__50214\,
            ce => \N__42640\,
            sr => \N__49632\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42763\,
            in1 => \N__42338\,
            in2 => \_gnd_net_\,
            in3 => \N__42322\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__50214\,
            ce => \N__42640\,
            sr => \N__49632\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42760\,
            in1 => \N__42318\,
            in2 => \_gnd_net_\,
            in3 => \N__42304\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__50214\,
            ce => \N__42640\,
            sr => \N__49632\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__42654\,
            in1 => \N__42761\,
            in2 => \_gnd_net_\,
            in3 => \N__42658\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50214\,
            ce => \N__42640\,
            sr => \N__49632\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42601\,
            in2 => \N__45390\,
            in3 => \N__45386\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47356\,
            in2 => \_gnd_net_\,
            in3 => \N__42580\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46825\,
            in2 => \_gnd_net_\,
            in3 => \N__42565\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47344\,
            in2 => \_gnd_net_\,
            in3 => \N__42562\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47338\,
            in2 => \_gnd_net_\,
            in3 => \N__42535\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47350\,
            in2 => \_gnd_net_\,
            in3 => \N__42532\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47362\,
            in2 => \_gnd_net_\,
            in3 => \N__42529\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47287\,
            in2 => \_gnd_net_\,
            in3 => \N__42973\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47320\,
            in2 => \_gnd_net_\,
            in3 => \N__42943\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47533\,
            in2 => \_gnd_net_\,
            in3 => \N__42913\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47332\,
            in2 => \_gnd_net_\,
            in3 => \N__42910\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47527\,
            in2 => \_gnd_net_\,
            in3 => \N__42883\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47326\,
            in2 => \_gnd_net_\,
            in3 => \N__42853\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47551\,
            in2 => \_gnd_net_\,
            in3 => \N__42823\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47371\,
            in3 => \N__42793\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47545\,
            in2 => \_gnd_net_\,
            in3 => \N__42790\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43399\,
            in2 => \_gnd_net_\,
            in3 => \N__43138\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43177\,
            in2 => \_gnd_net_\,
            in3 => \N__43135\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43342\,
            in2 => \_gnd_net_\,
            in3 => \N__43114\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43384\,
            in2 => \_gnd_net_\,
            in3 => \N__43093\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43417\,
            in2 => \_gnd_net_\,
            in3 => \N__43063\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43408\,
            in2 => \_gnd_net_\,
            in3 => \N__43030\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47539\,
            in2 => \_gnd_net_\,
            in3 => \N__43027\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43333\,
            in2 => \_gnd_net_\,
            in3 => \N__43003\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43390\,
            in2 => \_gnd_net_\,
            in3 => \N__43291\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43726\,
            in2 => \_gnd_net_\,
            in3 => \N__43258\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44281\,
            in3 => \N__43255\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43717\,
            in3 => \N__43228\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43672\,
            in2 => \_gnd_net_\,
            in3 => \N__43204\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43201\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43189\,
            in3 => \N__46801\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48049\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46803\,
            in1 => \N__48529\,
            in2 => \N__46418\,
            in3 => \N__43170\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47926\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48559\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48085\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48451\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47967\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48086\,
            in1 => \N__46802\,
            in2 => \N__46419\,
            in3 => \N__43371\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48005\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48485\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48373\,
            in1 => \N__46819\,
            in2 => \N__46420\,
            in3 => \N__43320\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48403\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48326\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__46818\,
            in1 => \N__43701\,
            in2 => \N__46379\,
            in3 => \N__48455\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48284\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_17_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43663\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44178\,
            in2 => \_gnd_net_\,
            in3 => \N__43452\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__43616\,
            in1 => \N__43590\,
            in2 => \N__43540\,
            in3 => \N__43537\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111001111"
        )
    port map (
            in0 => \N__45122\,
            in1 => \N__45297\,
            in2 => \N__44832\,
            in3 => \N__43486\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \N__49611\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000110101111"
        )
    port map (
            in0 => \N__45296\,
            in1 => \N__45123\,
            in2 => \N__44833\,
            in3 => \N__43429\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \N__49611\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIKOBP_17_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44265\,
            in1 => \N__44081\,
            in2 => \N__44140\,
            in3 => \N__44236\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIKOBPZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43785\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44179\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44135\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI898P_14_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44080\,
            in1 => \N__43872\,
            in2 => \N__43793\,
            in3 => \N__43837\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI898PZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45118\,
            in1 => \N__45309\,
            in2 => \N__44806\,
            in3 => \N__43813\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50248\,
            ce => 'H',
            sr => \N__49615\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011111110"
        )
    port map (
            in0 => \N__45307\,
            in1 => \N__45120\,
            in2 => \N__44808\,
            in3 => \N__43750\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50248\,
            ce => 'H',
            sr => \N__49615\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__45119\,
            in1 => \N__45310\,
            in2 => \N__44807\,
            in3 => \N__43738\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50248\,
            ce => 'H',
            sr => \N__49615\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011111110"
        )
    port map (
            in0 => \N__45308\,
            in1 => \N__45121\,
            in2 => \N__44809\,
            in3 => \N__44947\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50248\,
            ce => 'H',
            sr => \N__49615\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44625\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44577\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44489\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44431\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2P9P1_20_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44395\,
            in1 => \N__44383\,
            in2 => \N__44371\,
            in3 => \N__44356\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44331\,
            lcout => \delay_measurement_inst.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50236\,
            ce => \N__49815\,
            sr => \N__49619\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48374\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46756\,
            in1 => \N__47448\,
            in2 => \N__46423\,
            in3 => \N__45570\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47863\,
            in1 => \N__46757\,
            in2 => \N__46421\,
            in3 => \N__47080\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46758\,
            in1 => \N__48143\,
            in2 => \N__46422\,
            in3 => \N__45516\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47862\,
            in1 => \N__47215\,
            in2 => \_gnd_net_\,
            in3 => \N__47079\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_1_25_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46798\,
            in2 => \_gnd_net_\,
            in3 => \N__46339\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__47219\,
            in1 => \N__48057\,
            in2 => \_gnd_net_\,
            in3 => \N__45440\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47300\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__47301\,
            in1 => \_gnd_net_\,
            in2 => \N__45367\,
            in3 => \N__47188\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48845\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50224\,
            ce => \N__48268\,
            sr => \N__49627\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48814\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50224\,
            ce => \N__48268\,
            sr => \N__49627\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47785\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__47192\,
            in1 => \N__47136\,
            in2 => \_gnd_net_\,
            in3 => \N__47508\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46706\,
            in1 => \N__47674\,
            in2 => \N__46408\,
            in3 => \N__47112\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46705\,
            in1 => \N__47861\,
            in2 => \N__46407\,
            in3 => \N__47078\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__47050\,
            in1 => \N__47035\,
            in2 => \_gnd_net_\,
            in3 => \N__46965\,
            lcout => \current_shift_inst.control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47011\,
            in2 => \N__46991\,
            in3 => \N__46849\,
            lcout => \current_shift_inst.control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47469\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46796\,
            in1 => \N__47822\,
            in2 => \N__46406\,
            in3 => \N__47400\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48175\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47821\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47507\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47860\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47437\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47893\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47665\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47578\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47732\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48220\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48133\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48530\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47701\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47620\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48741\,
            in2 => \N__48810\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__50195\,
            ce => \N__48266\,
            sr => \N__49651\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48717\,
            in2 => \N__48774\,
            in3 => \N__47452\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__50195\,
            ce => \N__48266\,
            sr => \N__49651\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48742\,
            in2 => \N__48696\,
            in3 => \N__47410\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__50195\,
            ce => \N__48266\,
            sr => \N__49651\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48718\,
            in2 => \N__48670\,
            in3 => \N__47866\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__50195\,
            ce => \N__48266\,
            sr => \N__49651\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48636\,
            in2 => \N__48697\,
            in3 => \N__47836\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__50195\,
            ce => \N__48266\,
            sr => \N__49651\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48666\,
            in2 => \N__48615\,
            in3 => \N__47803\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__50195\,
            ce => \N__48266\,
            sr => \N__49651\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48637\,
            in2 => \N__49066\,
            in3 => \N__47758\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__50195\,
            ce => \N__48266\,
            sr => \N__49651\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49038\,
            in2 => \N__48616\,
            in3 => \N__47716\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__50195\,
            ce => \N__48266\,
            sr => \N__49651\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49065\,
            in2 => \N__49014\,
            in3 => \N__47677\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__50188\,
            ce => \N__48265\,
            sr => \N__49655\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49039\,
            in2 => \N__48987\,
            in3 => \N__47638\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__50188\,
            ce => \N__48265\,
            sr => \N__49655\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48960\,
            in2 => \N__49015\,
            in3 => \N__47593\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__50188\,
            ce => \N__48265\,
            sr => \N__49655\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48933\,
            in2 => \N__48988\,
            in3 => \N__47554\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__50188\,
            ce => \N__48265\,
            sr => \N__49655\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48961\,
            in2 => \N__48906\,
            in3 => \N__48193\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__50188\,
            ce => \N__48265\,
            sr => \N__49655\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48876\,
            in2 => \N__48937\,
            in3 => \N__48148\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__50188\,
            ce => \N__48265\,
            sr => \N__49655\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49311\,
            in2 => \N__48907\,
            in3 => \N__48103\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__50188\,
            ce => \N__48265\,
            sr => \N__49655\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48877\,
            in2 => \N__49285\,
            in3 => \N__48067\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__50188\,
            ce => \N__48265\,
            sr => \N__49655\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49312\,
            in2 => \N__49254\,
            in3 => \N__48022\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__50182\,
            ce => \N__48263\,
            sr => \N__49661\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49284\,
            in2 => \N__49224\,
            in3 => \N__47989\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__50182\,
            ce => \N__48263\,
            sr => \N__49661\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49194\,
            in2 => \N__49255\,
            in3 => \N__47956\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__50182\,
            ce => \N__48263\,
            sr => \N__49661\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49170\,
            in2 => \N__49225\,
            in3 => \N__47908\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__50182\,
            ce => \N__48263\,
            sr => \N__49661\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49195\,
            in2 => \N__49146\,
            in3 => \N__48541\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__50182\,
            ce => \N__48263\,
            sr => \N__49661\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49171\,
            in2 => \N__49119\,
            in3 => \N__48505\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__50182\,
            ce => \N__48263\,
            sr => \N__49661\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49092\,
            in2 => \N__49147\,
            in3 => \N__48469\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__50182\,
            ce => \N__48263\,
            sr => \N__49661\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50631\,
            in2 => \N__49120\,
            in3 => \N__48430\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__50182\,
            ce => \N__48263\,
            sr => \N__49661\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49093\,
            in2 => \N__50604\,
            in3 => \N__48385\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_18_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__50177\,
            ce => \N__48262\,
            sr => \N__49666\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50632\,
            in2 => \N__50577\,
            in3 => \N__48346\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__50177\,
            ce => \N__48262\,
            sr => \N__49666\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50551\,
            in2 => \N__50605\,
            in3 => \N__48310\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__50177\,
            ce => \N__48262\,
            sr => \N__49666\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50407\,
            in2 => \N__50578\,
            in3 => \N__48271\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__50177\,
            ce => \N__48262\,
            sr => \N__49666\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48238\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50520\,
            in1 => \N__48797\,
            in2 => \_gnd_net_\,
            in3 => \N__48781\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_22_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__50172\,
            ce => \N__50389\,
            sr => \N__49673\
        );

    \current_shift_inst.timer_s1.counter_1_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50504\,
            in1 => \N__48764\,
            in2 => \_gnd_net_\,
            in3 => \N__48745\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__50172\,
            ce => \N__50389\,
            sr => \N__49673\
        );

    \current_shift_inst.timer_s1.counter_2_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50521\,
            in1 => \N__48735\,
            in2 => \_gnd_net_\,
            in3 => \N__48721\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__50172\,
            ce => \N__50389\,
            sr => \N__49673\
        );

    \current_shift_inst.timer_s1.counter_3_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50505\,
            in1 => \N__48716\,
            in2 => \_gnd_net_\,
            in3 => \N__48700\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__50172\,
            ce => \N__50389\,
            sr => \N__49673\
        );

    \current_shift_inst.timer_s1.counter_4_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50522\,
            in1 => \N__48689\,
            in2 => \_gnd_net_\,
            in3 => \N__48673\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__50172\,
            ce => \N__50389\,
            sr => \N__49673\
        );

    \current_shift_inst.timer_s1.counter_5_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50506\,
            in1 => \N__48662\,
            in2 => \_gnd_net_\,
            in3 => \N__48640\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__50172\,
            ce => \N__50389\,
            sr => \N__49673\
        );

    \current_shift_inst.timer_s1.counter_6_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50523\,
            in1 => \N__48635\,
            in2 => \_gnd_net_\,
            in3 => \N__48619\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__50172\,
            ce => \N__50389\,
            sr => \N__49673\
        );

    \current_shift_inst.timer_s1.counter_7_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50507\,
            in1 => \N__48603\,
            in2 => \_gnd_net_\,
            in3 => \N__48589\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__50172\,
            ce => \N__50389\,
            sr => \N__49673\
        );

    \current_shift_inst.timer_s1.counter_8_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50511\,
            in1 => \N__49061\,
            in2 => \_gnd_net_\,
            in3 => \N__49042\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_23_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__50166\,
            ce => \N__50385\,
            sr => \N__49680\
        );

    \current_shift_inst.timer_s1.counter_9_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50515\,
            in1 => \N__49037\,
            in2 => \_gnd_net_\,
            in3 => \N__49018\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__50166\,
            ce => \N__50385\,
            sr => \N__49680\
        );

    \current_shift_inst.timer_s1.counter_10_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50508\,
            in1 => \N__49007\,
            in2 => \_gnd_net_\,
            in3 => \N__48991\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__50166\,
            ce => \N__50385\,
            sr => \N__49680\
        );

    \current_shift_inst.timer_s1.counter_11_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50512\,
            in1 => \N__48980\,
            in2 => \_gnd_net_\,
            in3 => \N__48964\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__50166\,
            ce => \N__50385\,
            sr => \N__49680\
        );

    \current_shift_inst.timer_s1.counter_12_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50509\,
            in1 => \N__48954\,
            in2 => \_gnd_net_\,
            in3 => \N__48940\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__50166\,
            ce => \N__50385\,
            sr => \N__49680\
        );

    \current_shift_inst.timer_s1.counter_13_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50513\,
            in1 => \N__48926\,
            in2 => \_gnd_net_\,
            in3 => \N__48910\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__50166\,
            ce => \N__50385\,
            sr => \N__49680\
        );

    \current_shift_inst.timer_s1.counter_14_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50510\,
            in1 => \N__48894\,
            in2 => \_gnd_net_\,
            in3 => \N__48880\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__50166\,
            ce => \N__50385\,
            sr => \N__49680\
        );

    \current_shift_inst.timer_s1.counter_15_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50514\,
            in1 => \N__48875\,
            in2 => \_gnd_net_\,
            in3 => \N__48859\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__50166\,
            ce => \N__50385\,
            sr => \N__49680\
        );

    \current_shift_inst.timer_s1.counter_16_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50524\,
            in1 => \N__49304\,
            in2 => \_gnd_net_\,
            in3 => \N__49288\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_18_24_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__50162\,
            ce => \N__50384\,
            sr => \N__49687\
        );

    \current_shift_inst.timer_s1.counter_17_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50516\,
            in1 => \N__49274\,
            in2 => \_gnd_net_\,
            in3 => \N__49258\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__50162\,
            ce => \N__50384\,
            sr => \N__49687\
        );

    \current_shift_inst.timer_s1.counter_18_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50525\,
            in1 => \N__49242\,
            in2 => \_gnd_net_\,
            in3 => \N__49228\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__50162\,
            ce => \N__50384\,
            sr => \N__49687\
        );

    \current_shift_inst.timer_s1.counter_19_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50517\,
            in1 => \N__49212\,
            in2 => \_gnd_net_\,
            in3 => \N__49198\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__50162\,
            ce => \N__50384\,
            sr => \N__49687\
        );

    \current_shift_inst.timer_s1.counter_20_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50526\,
            in1 => \N__49188\,
            in2 => \_gnd_net_\,
            in3 => \N__49174\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__50162\,
            ce => \N__50384\,
            sr => \N__49687\
        );

    \current_shift_inst.timer_s1.counter_21_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50518\,
            in1 => \N__49164\,
            in2 => \_gnd_net_\,
            in3 => \N__49150\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__50162\,
            ce => \N__50384\,
            sr => \N__49687\
        );

    \current_shift_inst.timer_s1.counter_22_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50527\,
            in1 => \N__49139\,
            in2 => \_gnd_net_\,
            in3 => \N__49123\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__50162\,
            ce => \N__50384\,
            sr => \N__49687\
        );

    \current_shift_inst.timer_s1.counter_23_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50519\,
            in1 => \N__49112\,
            in2 => \_gnd_net_\,
            in3 => \N__49096\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__50162\,
            ce => \N__50384\,
            sr => \N__49687\
        );

    \current_shift_inst.timer_s1.counter_24_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50528\,
            in1 => \N__49085\,
            in2 => \_gnd_net_\,
            in3 => \N__49069\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_18_25_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__50159\,
            ce => \N__50383\,
            sr => \N__49692\
        );

    \current_shift_inst.timer_s1.counter_25_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50532\,
            in1 => \N__50624\,
            in2 => \_gnd_net_\,
            in3 => \N__50608\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__50159\,
            ce => \N__50383\,
            sr => \N__49692\
        );

    \current_shift_inst.timer_s1.counter_26_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50529\,
            in1 => \N__50597\,
            in2 => \_gnd_net_\,
            in3 => \N__50581\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__50159\,
            ce => \N__50383\,
            sr => \N__49692\
        );

    \current_shift_inst.timer_s1.counter_27_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50533\,
            in1 => \N__50570\,
            in2 => \_gnd_net_\,
            in3 => \N__50554\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__50159\,
            ce => \N__50383\,
            sr => \N__49692\
        );

    \current_shift_inst.timer_s1.counter_28_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50530\,
            in1 => \N__50550\,
            in2 => \_gnd_net_\,
            in3 => \N__50536\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__50159\,
            ce => \N__50383\,
            sr => \N__49692\
        );

    \current_shift_inst.timer_s1.counter_29_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__50403\,
            in1 => \N__50531\,
            in2 => \_gnd_net_\,
            in3 => \N__50410\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50159\,
            ce => \N__50383\,
            sr => \N__49692\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50332\,
            lcout => \delay_measurement_inst.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50249\,
            ce => \N__49816\,
            sr => \N__49620\
        );
end \INTERFACE\;
